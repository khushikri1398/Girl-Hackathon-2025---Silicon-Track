
module simple_alu_0580(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0580
);

    always @(*) begin
        case(op)
            
            4'd0: result_0580 = (((b << 3) & (((14'd11019 ^ b) ? 14'd916 : 7170) * ((14'd12119 ? 14'd644 : 1452) + 14'd7097))) * ((((14'd207 >> 1) >> 2) + a) & (((14'd7424 & 14'd13938) ? a : 1736) ^ 14'd11565)));
            
            4'd1: result_0580 = (a + a);
            
            4'd2: result_0580 = ((~(((14'd11964 << 2) << 3) * (14'd6661 << 2))) * (((b >> 2) ^ 14'd11208) >> 1));
            
            4'd3: result_0580 = ((14'd6722 << 3) << 3);
            
            4'd4: result_0580 = ((~b) * 14'd2872);
            
            4'd5: result_0580 = (((~((14'd11484 | a) & (~b))) & (((14'd12850 & b) - (a + 14'd4191)) + ((14'd11648 << 3) & (a ? 14'd2436 : 7783)))) * ((14'd13589 | (b ^ 14'd3455)) << 1));
            
            4'd6: result_0580 = (b | ((((14'd1255 + 14'd7097) >> 1) >> 2) * (((14'd2726 - b) << 3) >> 3)));
            
            4'd7: result_0580 = ((14'd10614 >> 3) - ((a - ((14'd8151 >> 1) ? 14'd7830 : 3069)) + (((a >> 2) << 1) + a)));
            
            4'd8: result_0580 = (((((14'd11231 << 2) ^ (~14'd3401)) | (~(14'd8471 | 14'd5254))) * (((14'd15587 ^ 14'd14735) & 14'd1777) ? (b - 14'd5991) : 6658)) ? (((a & (14'd10416 & a)) - 14'd6062) >> 1) : 4752);
            
            4'd9: result_0580 = (((14'd6196 & (14'd1662 | (14'd1792 | a))) + b) & (14'd10147 | (((a | a) ? (14'd15967 << 1) : 5806) | ((14'd15309 & 14'd627) ? (b & 14'd7761) : 13447))));
            
            default: result_0580 = 14'd12754;
        endcase
    end

endmodule
        