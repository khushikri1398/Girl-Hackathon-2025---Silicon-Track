
module simple_alu_0479(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0479
);

    always @(*) begin
        case(op)
            
            4'd0: result_0479 = (((~a) + ((b + b) >> 3)) | b);
            
            4'd1: result_0479 = ((((12'd1542 ? a : 1960) >> 2) + 12'd3110) * ((~(a >> 1)) & ((12'd1122 & 12'd3870) & (a ? b : 2022))));
            
            4'd2: result_0479 = ((12'd1640 + ((~a) << 2)) | ((~b) | (a << 1)));
            
            4'd3: result_0479 = ((((12'd11 + a) & (b * b)) & ((a | a) >> 2)) - 12'd2260);
            
            4'd4: result_0479 = ((~b) ^ ((a | (12'd2388 << 1)) + b));
            
            4'd5: result_0479 = (a >> 3);
            
            4'd6: result_0479 = ((~((b | a) & (a - 12'd1255))) << 2);
            
            4'd7: result_0479 = (((12'd1586 << 1) & ((12'd3077 ? 12'd1254 : 724) | (a | a))) ^ b);
            
            4'd8: result_0479 = (a | (((a ^ 12'd796) + 12'd733) >> 3));
            
            4'd9: result_0479 = ((a + b) >> 3);
            
            4'd10: result_0479 = (((12'd66 | a) ^ 12'd3486) >> 3);
            
            4'd11: result_0479 = ((12'd3070 & ((b | b) ^ 12'd2435)) ? (((a ? a : 2975) ^ (a * b)) | (12'd4027 << 3)) : 1419);
            
            4'd12: result_0479 = (~12'd598);
            
            4'd13: result_0479 = (a - (((12'd661 * 12'd1349) - (a << 2)) - b));
            
            4'd14: result_0479 = ((b >> 3) + 12'd758);
            
            default: result_0479 = 12'd399;
        endcase
    end

endmodule
        