
module simple_alu_0125(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0125
);

    always @(*) begin
        case(op)
            
            4'd0: result_0125 = (14'd5128 ^ (a << 2));
            
            4'd1: result_0125 = (14'd3247 - b);
            
            4'd2: result_0125 = (14'd931 - ((((b - 14'd1882) >> 2) | ((a << 2) | (a - a))) >> 3));
            
            4'd3: result_0125 = ((((14'd11878 ? (14'd3695 ? 14'd6680 : 3256) : 5794) - (14'd10738 << 2)) ? (((14'd7178 + b) - a) >> 3) : 12914) >> 2);
            
            4'd4: result_0125 = (14'd9354 ? 14'd2464 : 6952);
            
            4'd5: result_0125 = (14'd7346 | 14'd16176);
            
            4'd6: result_0125 = (a | (~(((b & 14'd15394) ? 14'd5487 : 8569) * ((b | 14'd13754) >> 2))));
            
            4'd7: result_0125 = ((a & (~(~(14'd5289 * 14'd3698)))) << 2);
            
            4'd8: result_0125 = ((((a >> 2) & (14'd12386 ^ (14'd6508 + 14'd3592))) + (~14'd12531)) & (14'd2908 << 1));
            
            4'd9: result_0125 = ((a ^ (((14'd12481 << 3) >> 1) ? b : 2355)) ^ ((((b ^ a) * 14'd495) + ((14'd9208 + b) ^ (14'd6447 | 14'd15378))) << 2));
            
            4'd10: result_0125 = ((((a | 14'd6672) ^ (14'd5070 * 14'd3259)) >> 1) << 1);
            
            4'd11: result_0125 = ((b | (((14'd6803 ? b : 4328) << 2) ? ((14'd13423 ? a : 3992) | (a << 1)) : 16129)) ? a : 8895);
            
            4'd12: result_0125 = ((((a >> 2) ? 14'd2250 : 6340) ^ 14'd14797) << 2);
            
            4'd13: result_0125 = ((~14'd14663) << 3);
            
            4'd14: result_0125 = ((~(a + 14'd15340)) + ((14'd13576 * b) - (14'd8360 * ((b - 14'd13851) & 14'd14183))));
            
            4'd15: result_0125 = ((14'd10332 ^ 14'd5372) | ((14'd3375 | a) | (14'd3816 - a)));
            
            default: result_0125 = 14'd8783;
        endcase
    end

endmodule
        