
module simple_alu_0427(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0427
);

    always @(*) begin
        case(op)
            
            4'd0: result_0427 = (14'd979 ^ (((~(14'd4037 ? b : 1140)) >> 1) ? ((~14'd9699) & ((14'd16113 ^ 14'd12134) ^ (a | b))) : 4103));
            
            4'd1: result_0427 = (((b | ((b & 14'd6907) + 14'd8990)) << 3) ^ a);
            
            4'd2: result_0427 = (((14'd13113 ? (14'd15474 >> 1) : 11728) * a) - ((((a * 14'd10293) + 14'd540) ? 14'd3890 : 4242) >> 1));
            
            4'd3: result_0427 = (((14'd14631 | ((b ^ 14'd8872) - b)) | (((14'd2166 + 14'd14624) | (14'd8757 + 14'd1124)) >> 2)) + ((((b - 14'd9527) - (b + 14'd2736)) << 1) | b));
            
            4'd4: result_0427 = ((14'd5388 + (b | 14'd10538)) >> 2);
            
            4'd5: result_0427 = (14'd12334 ? ((((14'd302 << 2) >> 1) | (b | (14'd16124 | 14'd13802))) - (~(14'd11235 - (14'd10439 * 14'd13446)))) : 7190);
            
            4'd6: result_0427 = ((14'd14133 * ((~(14'd3317 & 14'd7900)) | ((a << 3) | (14'd4273 * a)))) * b);
            
            4'd7: result_0427 = ((14'd5221 ^ 14'd15227) ? (~(((14'd5076 | 14'd16280) - b) | a)) : 5627);
            
            4'd8: result_0427 = (((((14'd8260 ^ 14'd10203) ^ (a ? 14'd1477 : 6868)) + ((14'd2899 ^ 14'd10982) ^ (a + 14'd6699))) | (((14'd12733 + b) * a) >> 2)) * ((b >> 3) & (~14'd11816)));
            
            4'd9: result_0427 = (((~(14'd4977 | (14'd941 ^ 14'd12063))) << 2) + 14'd265);
            
            4'd10: result_0427 = ((((a * 14'd8878) ^ ((~14'd15918) * 14'd1094)) << 3) - ((((a >> 1) + (14'd9540 * 14'd6993)) << 1) - b));
            
            4'd11: result_0427 = (b - 14'd12868);
            
            4'd12: result_0427 = (((14'd2181 | ((a << 3) ^ b)) & 14'd5218) >> 2);
            
            4'd13: result_0427 = (~((((a & a) * (14'd12982 & a)) ? (14'd7510 + (14'd5550 + 14'd2819)) : 10612) * ((~(14'd573 & b)) + ((14'd15255 ? 14'd11002 : 4004) & (14'd1381 ^ a)))));
            
            default: result_0427 = a;
        endcase
    end

endmodule
        