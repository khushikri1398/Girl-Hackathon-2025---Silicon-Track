
module simple_alu_0028(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0028
);

    always @(*) begin
        case(op)
            
            4'd0: result_0028 = ((14'd11852 - (((~14'd8690) >> 1) | ((b ^ 14'd1479) | (b | 14'd13763)))) ^ (((b ? (b ? 14'd15758 : 10535) : 1921) + (14'd2032 & (14'd4387 | 14'd724))) >> 3));
            
            4'd1: result_0028 = (((14'd1135 >> 3) << 2) * ((((~14'd6627) + (14'd603 << 2)) + ((a ? a : 6985) * 14'd1150)) ? (~((a ? b : 5591) >> 2)) : 14729));
            
            4'd2: result_0028 = (((((14'd1867 | a) + (14'd3162 ^ 14'd2766)) ^ a) | 14'd13027) >> 1);
            
            4'd3: result_0028 = (((14'd5499 | ((14'd2175 & a) * (14'd13265 * a))) << 1) << 1);
            
            4'd4: result_0028 = (~(b ? (((b ^ a) ^ b) * ((14'd2929 ^ 14'd7310) + (b & a))) : 6425));
            
            4'd5: result_0028 = (b + ((((a | 14'd8830) & (b * 14'd1146)) | ((14'd8287 & 14'd10691) + (a - 14'd2399))) ^ ((~(14'd2692 ^ a)) | ((b << 1) & 14'd5272))));
            
            4'd6: result_0028 = (((b >> 3) >> 2) & ((((14'd3556 - a) >> 3) << 3) ? (b >> 1) : 1353));
            
            4'd7: result_0028 = ((14'd3912 ? (14'd10487 + a) : 7519) + 14'd7712);
            
            4'd8: result_0028 = (14'd4381 ? ((~((14'd3617 << 2) ? (b ? 14'd15363 : 12773) : 8686)) ? b : 603) : 16365);
            
            4'd9: result_0028 = (b >> 2);
            
            default: result_0028 = 14'd16329;
        endcase
    end

endmodule
        