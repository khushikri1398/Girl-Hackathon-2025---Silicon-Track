
module simple_alu_0817(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0817
);

    always @(*) begin
        case(op)
            
            4'd0: result_0817 = ((b * 14'd6093) * (~(((14'd4058 - 14'd1200) ^ (a + b)) & ((14'd2948 ^ 14'd6015) & 14'd15783))));
            
            4'd1: result_0817 = (a << 1);
            
            4'd2: result_0817 = (((((14'd14605 ^ b) & (14'd15586 >> 3)) >> 1) | (((b * a) << 3) << 2)) ? 14'd14875 : 3626);
            
            4'd3: result_0817 = (((a & b) ? (((b + 14'd4552) | (14'd9302 ^ a)) >> 1) : 4781) * (14'd15627 ? (((a | a) << 3) ^ ((a << 1) ^ (b * 14'd1408))) : 7567));
            
            4'd4: result_0817 = (a << 2);
            
            4'd5: result_0817 = (((((~14'd6051) ^ (a * 14'd4588)) * 14'd718) * (14'd6153 << 3)) - 14'd10285);
            
            4'd6: result_0817 = ((((14'd6742 * (b - 14'd1886)) >> 1) >> 2) - b);
            
            4'd7: result_0817 = (((((a | a) - 14'd7606) << 1) >> 3) & a);
            
            4'd8: result_0817 = (a ? (((b + (b >> 2)) & 14'd11991) >> 3) : 12256);
            
            4'd9: result_0817 = (((((b * 14'd2941) ^ (14'd758 | 14'd14826)) * 14'd7085) ? (~(a * (14'd8210 ^ 14'd15615))) : 8998) + ((((b << 1) * (14'd14081 - 14'd12612)) + (~(14'd13484 + a))) ? (((a + a) - (14'd5934 ^ a)) >> 3) : 5416));
            
            4'd10: result_0817 = (14'd9804 >> 2);
            
            4'd11: result_0817 = (~a);
            
            default: result_0817 = 14'd10577;
        endcase
    end

endmodule
        