
module simple_alu_0356(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0356
);

    always @(*) begin
        case(op)
            
            4'd0: result_0356 = ((14'd6915 ? (14'd4133 + ((14'd12701 ? 14'd7751 : 9158) + (a + b))) : 7254) - 14'd4045);
            
            4'd1: result_0356 = ((~((14'd5453 << 1) * ((14'd14514 | 14'd5014) | (~14'd4238)))) + (14'd2713 & (14'd3295 ^ a)));
            
            4'd2: result_0356 = (a - (((14'd9597 + (b & 14'd12588)) + 14'd10430) ^ 14'd6657));
            
            4'd3: result_0356 = (a | ((((14'd10517 & 14'd14977) << 1) | ((14'd7325 ? a : 6537) - 14'd7341)) - (14'd8413 << 2)));
            
            4'd4: result_0356 = (((((14'd9981 | 14'd5168) ? (14'd9597 ^ b) : 14985) >> 3) - 14'd5515) * 14'd5458);
            
            4'd5: result_0356 = (14'd5519 << 3);
            
            4'd6: result_0356 = ((~14'd9252) ^ (a ? 14'd3182 : 5381));
            
            4'd7: result_0356 = ((14'd12275 ^ (14'd1311 - ((14'd16003 >> 2) >> 3))) * (14'd11757 ? (a ? (14'd1746 * 14'd12595) : 13720) : 13154));
            
            4'd8: result_0356 = ((((14'd2378 & 14'd3047) - (14'd10143 >> 3)) ^ ((~(a + a)) >> 2)) & ((14'd10808 & ((a & 14'd8612) ? (b + b) : 14788)) << 3));
            
            4'd9: result_0356 = (~14'd15202);
            
            4'd10: result_0356 = (((((~14'd15933) >> 1) & ((~14'd9222) * b)) - (14'd2601 << 2)) - ((((14'd10151 & 14'd10994) + (a >> 2)) * (14'd10939 ? (a | 14'd6108) : 2811)) ? 14'd9514 : 9037));
            
            4'd11: result_0356 = (((b * (~14'd15793)) | b) * (((14'd5030 * (14'd13512 << 1)) + ((b << 2) & (14'd2241 * 14'd14169))) & (((14'd13911 << 2) + 14'd12003) >> 1)));
            
            4'd12: result_0356 = (14'd3847 * 14'd8679);
            
            4'd13: result_0356 = (((((b * b) ^ b) ? ((a ? 14'd3862 : 3856) + (~14'd7937)) : 7081) | 14'd3353) >> 2);
            
            4'd14: result_0356 = (14'd3773 | ((14'd7229 ^ a) * a));
            
            4'd15: result_0356 = (14'd8199 << 3);
            
            default: result_0356 = 14'd6485;
        endcase
    end

endmodule
        