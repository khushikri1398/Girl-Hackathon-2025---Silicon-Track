
module simple_alu_0786(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0786
);

    always @(*) begin
        case(op)
            
            4'd0: result_0786 = ((14'd16286 * (b * (~(14'd9659 + 14'd11385)))) >> 3);
            
            4'd1: result_0786 = ((14'd5337 >> 1) * (14'd14382 - (((14'd12088 << 2) << 3) >> 3)));
            
            4'd2: result_0786 = (~((((14'd10984 >> 2) ^ (14'd5045 >> 2)) >> 2) * (14'd4580 ? ((14'd7776 | 14'd14554) ^ 14'd6838) : 6129)));
            
            4'd3: result_0786 = ((~(((14'd7468 << 1) ? (14'd14201 - 14'd9561) : 3112) << 3)) >> 1);
            
            4'd4: result_0786 = (((b + (~(a >> 2))) ? ((~b) & 14'd2154) : 3651) ^ (((a - 14'd13065) - ((a - 14'd6906) ? 14'd2706 : 2846)) * ((~(14'd337 >> 3)) & ((14'd1191 | 14'd1394) << 2))));
            
            4'd5: result_0786 = (((a ? b : 15213) ^ (((14'd441 & b) >> 1) & (14'd7064 + (14'd11054 + a)))) | a);
            
            default: result_0786 = a;
        endcase
    end

endmodule
        