
module simple_alu_0736(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0736
);

    always @(*) begin
        case(op)
            
            4'd0: result_0736 = (14'd10402 >> 1);
            
            4'd1: result_0736 = ((~(((14'd1637 ? 14'd10487 : 7892) * (14'd14475 + 14'd14265)) | a)) ^ (((14'd6809 ? (~14'd5813) : 3106) >> 3) - (((b * 14'd6747) << 2) & 14'd10484)));
            
            4'd2: result_0736 = (a >> 1);
            
            4'd3: result_0736 = (((14'd10628 >> 1) | ((14'd15239 >> 2) >> 1)) | (((a << 2) | (a ^ (a & 14'd5527))) >> 3));
            
            4'd4: result_0736 = (((((a & 14'd413) + (b - 14'd5986)) & (a ^ (b & 14'd2572))) & a) + (a ^ (((b * b) + (~14'd5971)) | ((b * 14'd11916) | (14'd1328 & 14'd16099)))));
            
            4'd5: result_0736 = ((((14'd14524 * (14'd2014 ? 14'd12069 : 14115)) | b) ? a : 10037) << 3);
            
            4'd6: result_0736 = (14'd565 | 14'd12152);
            
            4'd7: result_0736 = ((a + (((a | a) << 3) + b)) >> 1);
            
            4'd8: result_0736 = (14'd1580 << 3);
            
            4'd9: result_0736 = ((~a) + ((((14'd8526 - b) ? b : 9266) ^ (14'd7223 & (14'd12549 ? b : 4623))) >> 1));
            
            4'd10: result_0736 = (((14'd6335 ? ((a * 14'd9710) ^ 14'd15166) : 2527) << 3) & 14'd4181);
            
            default: result_0736 = a;
        endcase
    end

endmodule
        