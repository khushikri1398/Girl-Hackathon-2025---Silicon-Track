
module simple_alu_0373(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0373
);

    always @(*) begin
        case(op)
            
            4'd0: result_0373 = (((b * b) & (a | ((a | 14'd1044) >> 3))) ^ 14'd4333);
            
            4'd1: result_0373 = (((14'd13953 ? b : 11744) & a) << 3);
            
            4'd2: result_0373 = (b << 1);
            
            4'd3: result_0373 = (~(~14'd11831));
            
            4'd4: result_0373 = ((14'd14437 - (((14'd2085 + a) * (a + a)) | b)) << 3);
            
            4'd5: result_0373 = (b * 14'd4075);
            
            4'd6: result_0373 = (((~(~(14'd15705 & 14'd8487))) & 14'd15951) | ((((b & 14'd7426) | (14'd5050 ? 14'd9046 : 16137)) << 1) | ((14'd12998 ^ (14'd244 ^ 14'd11956)) ? ((b * 14'd5399) >> 1) : 946)));
            
            4'd7: result_0373 = (((((14'd3394 >> 3) | 14'd13580) << 1) << 1) * (14'd3442 * (a >> 1)));
            
            4'd8: result_0373 = (((((a | b) >> 3) >> 2) & (((14'd11424 | 14'd765) ? (~14'd6336) : 15278) & ((14'd5 ? b : 3720) << 2))) - (((14'd2169 - (14'd7402 ^ b)) >> 3) ? (14'd10408 * ((a >> 1) + (~14'd11974))) : 6287));
            
            default: result_0373 = 14'd709;
        endcase
    end

endmodule
        