
module simple_alu_0662(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0662
);

    always @(*) begin
        case(op)
            
            4'd0: result_0662 = (a >> 3);
            
            4'd1: result_0662 = ((14'd9660 ? (((a + a) ? (14'd4471 << 1) : 301) >> 2) : 1865) ? ((14'd14630 - (b - (14'd15049 << 2))) * (((14'd1483 ? 14'd2335 : 15108) << 1) ? ((14'd14779 & a) >> 2) : 14575)) : 12106);
            
            4'd2: result_0662 = (a << 2);
            
            4'd3: result_0662 = ((~(14'd12241 ^ ((b << 3) << 2))) ^ ((14'd8283 | (~(14'd1886 + 14'd15711))) ^ (a * 14'd1771)));
            
            4'd4: result_0662 = (((14'd13675 << 1) >> 2) * ((a * 14'd4184) | 14'd3644));
            
            4'd5: result_0662 = ((((14'd510 - 14'd14302) - (~(14'd2714 >> 2))) & (((b >> 3) << 2) ? ((b ^ 14'd12247) - (~a)) : 960)) & 14'd946);
            
            4'd6: result_0662 = (14'd4374 | 14'd1259);
            
            4'd7: result_0662 = ((~(((a << 3) << 2) * (14'd13472 >> 1))) >> 3);
            
            4'd8: result_0662 = (14'd5868 ? (~14'd4400) : 14567);
            
            4'd9: result_0662 = ((14'd14664 | (((b >> 3) ? (b & 14'd4745) : 14138) & (14'd16038 ? (14'd9745 - 14'd9963) : 6079))) | 14'd461);
            
            4'd10: result_0662 = (((b << 2) | (((14'd11388 ^ a) & (b ? b : 14374)) & ((a * 14'd14724) & (14'd5614 >> 3)))) | ((((14'd9275 << 2) * (14'd14333 | b)) << 2) ^ (14'd14458 ? (14'd4110 | b) : 6923)));
            
            4'd11: result_0662 = ((a ^ (~(14'd11105 ^ (~b)))) & ((14'd13353 & 14'd4547) << 2));
            
            4'd12: result_0662 = (((((~14'd5308) - (14'd9032 * 14'd177)) >> 2) >> 3) ? ((((14'd3895 ? a : 14860) | (14'd15175 - 14'd9135)) * ((14'd3579 + 14'd10373) & (14'd2261 >> 1))) * (14'd6742 ^ ((14'd3879 ? 14'd13651 : 5567) ? (a | b) : 13780))) : 7906);
            
            4'd13: result_0662 = (14'd5474 >> 2);
            
            4'd14: result_0662 = (14'd6471 << 3);
            
            4'd15: result_0662 = ((14'd8300 + (~((14'd7458 << 2) * (14'd1676 + 14'd161)))) ^ b);
            
            default: result_0662 = b;
        endcase
    end

endmodule
        