
module simple_alu_0819(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0819
);

    always @(*) begin
        case(op)
            
            4'd0: result_0819 = (14'd4961 << 3);
            
            4'd1: result_0819 = (((~(~14'd2085)) | 14'd12202) >> 2);
            
            4'd2: result_0819 = (((14'd6842 + (~(b & 14'd13462))) | 14'd12036) | (~(((14'd4941 ? a : 10862) * (14'd14255 >> 2)) + 14'd15848)));
            
            4'd3: result_0819 = (a ? ((14'd6114 + ((14'd16109 * b) - 14'd14104)) - ((b & (b ? 14'd8043 : 14576)) - 14'd2545)) : 3725);
            
            4'd4: result_0819 = (14'd8405 + 14'd5776);
            
            4'd5: result_0819 = (((((14'd5379 + 14'd7710) | (14'd3529 | a)) * ((a - 14'd327) & (14'd15410 - a))) & (14'd5895 >> 2)) + (((14'd13001 << 1) * (~(a ? b : 5789))) + (((b * b) ? (14'd11978 << 3) : 5021) ^ ((14'd8048 ^ a) << 1))));
            
            4'd6: result_0819 = (((((b * 14'd2365) * (14'd13058 | 14'd2041)) ? (14'd10521 | (a | a)) : 12418) + (14'd12157 ? (14'd9821 >> 2) : 11654)) + ((((a ? 14'd984 : 14044) - (14'd7168 + b)) | b) ? (a & ((a >> 1) - (~14'd9516))) : 15993));
            
            4'd7: result_0819 = (((((14'd14005 ? b : 13359) ? (b * 14'd6318) : 2988) << 3) - (a >> 1)) | ((((14'd555 << 2) ? b : 9928) | a) | (((b * a) ? a : 4520) + ((b & 14'd8789) ^ (14'd13224 * a)))));
            
            4'd8: result_0819 = (14'd11140 * ((b >> 2) & (14'd4775 & a)));
            
            4'd9: result_0819 = (14'd3911 | 14'd15024);
            
            4'd10: result_0819 = ((~(~14'd11644)) << 2);
            
            4'd11: result_0819 = (((((b * 14'd14359) | (a + 14'd5515)) ^ (b << 3)) | (((14'd10728 ? b : 7442) & (a & 14'd10133)) << 1)) * (((~b) - ((b << 3) & 14'd3009)) ? (((a - 14'd3837) >> 1) | ((14'd3316 ? 14'd16169 : 6390) * (14'd10910 ^ a))) : 5518));
            
            4'd12: result_0819 = ((14'd4539 + (~(a ^ (14'd4651 >> 2)))) >> 1);
            
            4'd13: result_0819 = (((((b * 14'd11859) ^ (b * 14'd15104)) << 2) << 1) ^ (~b));
            
            4'd14: result_0819 = (14'd5428 >> 1);
            
            4'd15: result_0819 = ((((14'd12417 * 14'd2457) & ((14'd13075 - a) - (14'd6289 & 14'd5816))) >> 1) & a);
            
            default: result_0819 = 14'd5004;
        endcase
    end

endmodule
        