
module simple_alu_0459(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0459
);

    always @(*) begin
        case(op)
            
            4'd0: result_0459 = ((~14'd3572) - 14'd8369);
            
            4'd1: result_0459 = (((a * b) << 1) ? ((~(14'd15894 | 14'd1146)) - 14'd5317) : 1318);
            
            4'd2: result_0459 = (((~14'd3455) - ((14'd11076 & b) | ((14'd13322 & 14'd7721) >> 1))) - ((((14'd14545 << 1) >> 3) + 14'd13410) | (((14'd993 >> 2) | 14'd13685) ? 14'd3351 : 247)));
            
            4'd3: result_0459 = (((~((b + 14'd15889) >> 2)) >> 2) << 3);
            
            4'd4: result_0459 = (((((14'd12836 * b) ? (a >> 3) : 3338) - ((a | 14'd6479) | (~14'd4731))) ^ (~(~(14'd9367 >> 1)))) << 3);
            
            4'd5: result_0459 = ((~(b * a)) + ((14'd3499 ^ ((b << 1) << 3)) ^ b));
            
            4'd6: result_0459 = (14'd2015 ? ((14'd9937 >> 1) ^ (a & ((~a) - (~14'd8694)))) : 3895);
            
            4'd7: result_0459 = (~((((a ^ 14'd11511) << 3) & 14'd1570) ^ a));
            
            4'd8: result_0459 = (((14'd12576 + ((14'd4471 & a) * (14'd3728 - 14'd4048))) * 14'd13944) ^ 14'd15533);
            
            4'd9: result_0459 = (~14'd13869);
            
            4'd10: result_0459 = ((((b >> 1) ^ 14'd13819) | ((~14'd4032) ? (~(14'd9440 * b)) : 10922)) + (a >> 2));
            
            4'd11: result_0459 = (b * (b + (((14'd6314 << 1) & 14'd7294) & a)));
            
            default: result_0459 = 14'd6625;
        endcase
    end

endmodule
        