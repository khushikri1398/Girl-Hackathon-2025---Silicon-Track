
module simple_alu_0897(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0897
);

    always @(*) begin
        case(op)
            
            4'd0: result_0897 = ((((14'd3537 - (a | 14'd7855)) * ((b ^ b) << 2)) ^ (((b + 14'd9293) + (b * a)) - (a + b))) - ((~(b - (b | a))) & (((14'd3919 | 14'd8273) * 14'd7137) >> 2)));
            
            4'd1: result_0897 = (~((((b ^ b) & (14'd1812 + 14'd14986)) | ((a ? 14'd7500 : 12642) + 14'd3965)) << 1));
            
            4'd2: result_0897 = ((14'd8358 - ((14'd15066 >> 2) ^ ((a << 3) * (14'd7497 ^ 14'd7818)))) * ((((14'd10426 ? 14'd10333 : 2681) & b) & ((14'd13780 + 14'd7788) ^ (14'd16103 << 3))) >> 2));
            
            4'd3: result_0897 = (a ? 14'd5572 : 11251);
            
            4'd4: result_0897 = (~((((14'd7824 << 3) + (~a)) & 14'd14269) * ((14'd4301 + (b * 14'd8548)) & 14'd10878)));
            
            default: result_0897 = 14'd10960;
        endcase
    end

endmodule
        