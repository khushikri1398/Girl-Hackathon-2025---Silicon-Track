
module simple_alu_0445(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0445
);

    always @(*) begin
        case(op)
            
            4'd0: result_0445 = (14'd11408 & ((b << 1) + (b >> 3)));
            
            4'd1: result_0445 = ((((14'd12914 << 2) - ((14'd12178 * a) | a)) | (((14'd371 * a) - (a | 14'd8621)) - (14'd10103 & 14'd7662))) + b);
            
            4'd2: result_0445 = (a - a);
            
            4'd3: result_0445 = (b ? (~(((14'd3624 - 14'd15226) & (~14'd10905)) ^ 14'd11437)) : 12785);
            
            4'd4: result_0445 = ((~(~((14'd9774 | 14'd13893) * (14'd8155 & 14'd12183)))) << 3);
            
            4'd5: result_0445 = (((((a ? 14'd2076 : 8503) ? a : 13694) ? b : 4138) << 3) ^ (~14'd11889));
            
            4'd6: result_0445 = (((((14'd5869 * 14'd4308) - 14'd12298) >> 2) ^ (14'd14786 << 2)) * ((((a ^ 14'd6892) & (14'd3851 | a)) & (14'd14892 + (b >> 1))) >> 2));
            
            4'd7: result_0445 = (~((b << 1) << 1));
            
            4'd8: result_0445 = ((14'd8136 >> 3) ? 14'd10894 : 10898);
            
            4'd9: result_0445 = (14'd1117 ? ((~((14'd7230 & b) << 2)) ? (((~b) ^ (14'd7408 ? 14'd11478 : 1270)) * ((14'd13488 >> 3) ^ (b >> 1))) : 15761) : 15352);
            
            4'd10: result_0445 = (~((((~14'd48) * 14'd317) | ((14'd9158 - 14'd8060) & b)) >> 2));
            
            4'd11: result_0445 = ((14'd6951 & (((14'd1596 * 14'd4186) + (a << 2)) ^ (14'd5140 & 14'd2719))) - ((a ? (a & (14'd16278 ^ a)) : 569) ? ((14'd11525 & 14'd8057) & a) : 6594));
            
            default: result_0445 = 14'd8919;
        endcase
    end

endmodule
        