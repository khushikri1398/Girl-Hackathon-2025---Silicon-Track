
module simple_alu_0585(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0585
);

    always @(*) begin
        case(op)
            
            4'd0: result_0585 = (a >> 1);
            
            4'd1: result_0585 = (((b << 1) ? ((14'd10107 ? a : 7220) - 14'd311) : 15213) >> 2);
            
            4'd2: result_0585 = (b * ((((a - a) | (~b)) & ((14'd2763 * 14'd5026) + (a ? b : 986))) | 14'd2780));
            
            4'd3: result_0585 = (((((a * a) ? (b << 1) : 4148) ? b : 10562) * (((a + b) - (14'd11117 * 14'd12587)) & ((14'd8995 ^ 14'd3092) + a))) | (14'd15579 * (14'd5611 - 14'd1603)));
            
            4'd4: result_0585 = ((~a) | ((14'd6109 * ((14'd1514 | 14'd8386) | (b ? 14'd5701 : 2735))) | (((14'd5812 ^ a) ? (14'd8056 << 3) : 3293) - (14'd15087 * (14'd7179 ^ a)))));
            
            4'd5: result_0585 = ((b ? (b | ((14'd3476 & 14'd5115) | (14'd1576 ? 14'd4800 : 7219))) : 8438) + (14'd15025 << 2));
            
            4'd6: result_0585 = (b - ((~(14'd5094 | (14'd6271 | 14'd4389))) * (((14'd15522 * 14'd13209) << 2) >> 1)));
            
            4'd7: result_0585 = (((((a ^ a) - (14'd12186 ^ 14'd6577)) & (b * 14'd11057)) << 2) - (((14'd14806 << 3) ? ((14'd1804 & 14'd13776) ? b : 13637) : 7397) - 14'd15827));
            
            4'd8: result_0585 = ((a | (~14'd12916)) ? (((14'd8129 ^ 14'd14516) + a) + b) : 12387);
            
            4'd9: result_0585 = ((a >> 1) & ((((a << 2) + 14'd12334) >> 2) + (((b ^ a) & (14'd2323 & b)) | ((14'd4606 ^ 14'd588) - b))));
            
            4'd10: result_0585 = ((~(((14'd3381 - b) + (14'd11184 - 14'd4081)) | ((a ? 14'd1711 : 8240) | 14'd12581))) ^ (((14'd4719 | (14'd11427 | 14'd7924)) - b) - b));
            
            4'd11: result_0585 = (14'd14317 >> 1);
            
            4'd12: result_0585 = (~b);
            
            4'd13: result_0585 = (~((14'd13834 >> 1) | (((14'd3961 + 14'd2039) - (14'd2241 >> 3)) ? (a + (14'd11695 << 2)) : 11993)));
            
            4'd14: result_0585 = ((((14'd14132 & (14'd549 >> 3)) ? (14'd14347 ? (a & 14'd6940) : 2768) : 4027) - 14'd4258) >> 3);
            
            4'd15: result_0585 = (b ? b : 2676);
            
            default: result_0585 = b;
        endcase
    end

endmodule
        