
module simple_alu_0507(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0507
);

    always @(*) begin
        case(op)
            
            4'd0: result_0507 = (14'd9360 ^ 14'd11312);
            
            4'd1: result_0507 = (((((14'd8504 & 14'd8097) | b) + (14'd16334 << 3)) + 14'd4121) << 2);
            
            4'd2: result_0507 = (((b * (14'd4610 | (14'd4203 * b))) ^ 14'd5945) & ((14'd8237 << 1) << 3));
            
            4'd3: result_0507 = ((((14'd14457 << 3) * ((14'd4796 * 14'd2436) ^ b)) + ((14'd9308 | (~14'd12115)) - ((a - b) ? 14'd9575 : 6431))) * (((14'd63 - 14'd14590) << 1) - a));
            
            4'd4: result_0507 = (a + ((((14'd3173 - b) - (a >> 3)) * 14'd9465) ^ 14'd2756));
            
            4'd5: result_0507 = ((((~(a << 1)) & (14'd13295 + (~b))) ^ 14'd3511) + ((((a & a) | 14'd13759) ? a : 11098) | (a + ((a + 14'd14645) * (14'd587 | 14'd9271)))));
            
            4'd6: result_0507 = ((((~14'd12517) + ((a - a) - (~b))) + ((b - (a - 14'd610)) * ((b ? b : 6860) + (14'd3440 << 2)))) >> 3);
            
            4'd7: result_0507 = (((((a - a) * 14'd16289) - 14'd7774) - (14'd15609 + ((b ? 14'd9572 : 6874) + (~b)))) ? ((((14'd5075 * 14'd4763) ? a : 1069) >> 1) | (b ? 14'd15309 : 11359)) : 12631);
            
            4'd8: result_0507 = (((((b ? a : 12681) << 1) ^ 14'd16093) - (((14'd11308 + 14'd12636) ^ (14'd8178 + a)) << 1)) >> 2);
            
            4'd9: result_0507 = (((((a * a) | (14'd448 | 14'd8356)) - ((14'd6156 * 14'd16058) << 3)) & (((14'd6981 - a) << 2) | 14'd2540)) * 14'd6023);
            
            4'd10: result_0507 = (((~14'd2486) * (((~14'd10926) + (~14'd4941)) & ((b >> 3) | (~14'd2751)))) >> 1);
            
            4'd11: result_0507 = (((~((a | 14'd7650) | (14'd11005 ? b : 8760))) & (b * ((14'd2100 ? a : 10212) | (b ? 14'd9371 : 8328)))) ? (14'd3273 & (14'd10100 ? (~(b - 14'd9716)) : 3056)) : 10962);
            
            4'd12: result_0507 = (~((((14'd16134 * 14'd6596) << 1) | ((14'd7979 | 14'd5171) * (~14'd13951))) + (((a >> 2) + (b ^ a)) << 3)));
            
            4'd13: result_0507 = (((14'd3620 ^ a) & (((14'd7037 * a) >> 3) | (14'd11771 >> 2))) | ((b & (a & 14'd8337)) | ((a & a) * ((14'd7777 | 14'd5504) << 3))));
            
            default: result_0507 = 14'd2064;
        endcase
    end

endmodule
        