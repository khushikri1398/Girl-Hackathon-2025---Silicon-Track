
module simple_alu_0781(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0781
);

    always @(*) begin
        case(op)
            
            4'd0: result_0781 = (~(~14'd10669));
            
            4'd1: result_0781 = (a >> 1);
            
            4'd2: result_0781 = (((((14'd7563 ^ a) & (b - 14'd6659)) ? ((14'd12650 * 14'd7403) << 3) : 3814) - 14'd7426) & 14'd5002);
            
            4'd3: result_0781 = (a + (14'd15697 << 2));
            
            4'd4: result_0781 = (((((14'd9212 >> 1) ^ 14'd10497) + a) + (a ? ((14'd9656 * 14'd2539) ? 14'd11808 : 4399) : 7539)) & 14'd11233);
            
            4'd5: result_0781 = ((14'd10962 | (((b << 2) & (14'd9750 << 1)) >> 2)) - (14'd5987 ^ (14'd15092 ? ((14'd2251 * a) * (14'd14160 * b)) : 6254)));
            
            4'd6: result_0781 = ((((b ^ (a - a)) >> 2) ^ ((14'd1744 & (a ^ 14'd15489)) ^ ((14'd350 ? a : 896) & (b * a)))) - ((14'd4886 | ((14'd15258 ? a : 13200) & (b >> 2))) << 1));
            
            4'd7: result_0781 = (((~((14'd15257 ? b : 7083) << 2)) & b) & ((((14'd2015 * a) + (14'd3797 << 2)) & ((b & a) * 14'd13939)) << 1));
            
            4'd8: result_0781 = (14'd5350 >> 1);
            
            4'd9: result_0781 = (((b * ((14'd7193 - a) << 1)) * (b & ((14'd10426 ? b : 14649) * (14'd13764 << 3)))) & (~(((a - 14'd854) ? (14'd7154 + a) : 7462) ? ((14'd5611 * 14'd3833) | (b & a)) : 15398)));
            
            4'd10: result_0781 = (b | ((((b & 14'd10015) - (b ^ 14'd1557)) + (a >> 2)) & (~((14'd11084 * 14'd4643) ? 14'd7371 : 6798))));
            
            4'd11: result_0781 = ((((a * (14'd2367 | b)) + ((a * 14'd9842) ? 14'd8426 : 4110)) ^ (((14'd13863 & b) + (~14'd10413)) ^ b)) | a);
            
            4'd12: result_0781 = ((14'd9332 >> 3) & ((14'd1194 & (~a)) - 14'd11532));
            
            4'd13: result_0781 = ((14'd6016 & 14'd7188) - ((((b * 14'd15930) + (14'd15434 >> 1)) >> 3) >> 2));
            
            default: result_0781 = 14'd4518;
        endcase
    end

endmodule
        