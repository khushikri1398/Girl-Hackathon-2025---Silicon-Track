
module simple_alu_0472(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0472
);

    always @(*) begin
        case(op)
            
            4'd0: result_0472 = ((14'd4518 & (14'd12224 >> 1)) >> 1);
            
            4'd1: result_0472 = (((((a + 14'd12419) & 14'd6648) << 2) << 1) << 1);
            
            4'd2: result_0472 = (~(14'd12706 ? b : 13250));
            
            4'd3: result_0472 = (~(((a | 14'd895) >> 2) ? ((a ? b : 6089) >> 3) : 8831));
            
            4'd4: result_0472 = (((14'd15014 - 14'd16217) - ((~(b << 1)) ? (14'd3061 + b) : 1008)) ^ b);
            
            4'd5: result_0472 = (~((((14'd8572 * a) ^ (a << 1)) ^ (14'd3158 & (14'd8159 ? 14'd6305 : 2636))) ^ 14'd976));
            
            4'd6: result_0472 = (b >> 3);
            
            4'd7: result_0472 = (~(14'd6369 * (14'd4594 - (a * b))));
            
            4'd8: result_0472 = (b - b);
            
            4'd9: result_0472 = (((14'd12192 * ((b >> 3) | b)) - 14'd11775) << 2);
            
            4'd10: result_0472 = (((14'd11267 | a) ^ (((14'd14945 - a) - (14'd11636 | b)) ? ((14'd6726 ^ b) << 1) : 13702)) >> 1);
            
            4'd11: result_0472 = (~14'd8583);
            
            4'd12: result_0472 = ((14'd1029 ? (((~a) - (14'd9947 - 14'd13340)) - 14'd8749) : 2366) >> 3);
            
            4'd13: result_0472 = (14'd7111 << 1);
            
            default: result_0472 = b;
        endcase
    end

endmodule
        