
module simple_alu_0613(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0613
);

    always @(*) begin
        case(op)
            
            4'd0: result_0613 = ((b ^ (~((a * 14'd7958) - 14'd8583))) | ((~14'd6409) | (~(b ? (a + 14'd12928) : 11204))));
            
            4'd1: result_0613 = ((~((14'd7771 & (14'd12538 + 14'd9319)) ^ (~(14'd5910 & 14'd14092)))) ? a : 74);
            
            4'd2: result_0613 = (~((((14'd391 - 14'd3783) ? b : 1203) ? ((~14'd147) >> 3) : 6509) * (a * (14'd13144 + 14'd3219))));
            
            4'd3: result_0613 = ((a >> 3) ^ ((14'd9042 & ((14'd3003 + b) ^ (a ^ a))) - ((a & (b + 14'd10096)) + (14'd4945 ^ (b ^ 14'd6421)))));
            
            4'd4: result_0613 = ((~(((14'd7205 - 14'd11848) ? (14'd7290 | a) : 8059) & ((a >> 1) * 14'd11676))) * ((~((14'd12577 + 14'd15125) - (~b))) & (~14'd9333)));
            
            4'd5: result_0613 = (((14'd3121 - ((14'd1142 ^ 14'd2335) - (b ? b : 3805))) & (((~14'd1555) ? (a ? b : 5583) : 2450) + ((14'd16042 - a) ^ 14'd7660))) & ((((14'd823 << 2) + (a ^ 14'd319)) ^ ((14'd7591 + 14'd3494) ^ (b >> 3))) >> 2));
            
            4'd6: result_0613 = (14'd11469 * (14'd6905 - (14'd4586 << 1)));
            
            4'd7: result_0613 = ((((~(a ^ a)) >> 1) + (((14'd15389 << 1) - (14'd9814 * 14'd4657)) | a)) | (~(b >> 1)));
            
            4'd8: result_0613 = (a ^ 14'd1866);
            
            4'd9: result_0613 = (14'd3790 | (~(((14'd12752 - 14'd10689) + 14'd6568) - ((a >> 1) ? (b * 14'd588) : 12544))));
            
            4'd10: result_0613 = ((~14'd4666) ? ((((14'd11544 << 3) & 14'd8952) + 14'd11732) + (((14'd7319 & 14'd8242) | (14'd4953 - 14'd2525)) * a)) : 2362);
            
            4'd11: result_0613 = (14'd151 << 2);
            
            4'd12: result_0613 = (((a + ((14'd3850 << 1) | (b - a))) - a) >> 3);
            
            4'd13: result_0613 = (((((14'd8249 >> 1) * 14'd8809) << 2) & ((a * (14'd11335 ^ 14'd14323)) * 14'd129)) - (14'd13585 ? (14'd2123 << 1) : 11403));
            
            4'd14: result_0613 = (~((14'd1415 * (a | (~b))) ^ 14'd12941));
            
            4'd15: result_0613 = (~((((~14'd7155) >> 3) ? 14'd9485 : 926) >> 2));
            
            default: result_0613 = 14'd15714;
        endcase
    end

endmodule
        