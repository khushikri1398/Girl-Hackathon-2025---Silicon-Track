
module simple_alu_0490(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0490
);

    always @(*) begin
        case(op)
            
            4'd0: result_0490 = (((((14'd11028 << 3) + (~14'd15851)) << 1) >> 2) & (14'd7261 & ((14'd10052 ? (~a) : 8050) ? (b * 14'd312) : 1457)));
            
            4'd1: result_0490 = (((((~14'd15874) + (14'd3179 >> 3)) >> 3) * (((b ? 14'd4494 : 5304) & b) << 1)) * (14'd11347 << 3));
            
            4'd2: result_0490 = (b & (~((a ? b : 7241) + 14'd13468)));
            
            4'd3: result_0490 = (((((14'd15734 ^ 14'd9809) + (14'd398 << 2)) << 1) ? b : 11303) ? ((((b * a) << 2) + ((14'd518 >> 1) ^ 14'd14591)) * ((14'd4449 & (b - 14'd1354)) ? ((b & a) ^ 14'd13576) : 12933)) : 7655);
            
            4'd4: result_0490 = ((a >> 2) + ((a >> 3) >> 3));
            
            4'd5: result_0490 = (((b + ((b >> 3) + (14'd11257 ? 14'd5768 : 14625))) ? (((a + 14'd4836) & (14'd10145 | 14'd7645)) + ((a ^ a) << 2)) : 9840) & b);
            
            4'd6: result_0490 = ((a ? 14'd6957 : 1115) ^ (~((14'd5923 | (~14'd5546)) | b)));
            
            4'd7: result_0490 = (14'd9299 << 3);
            
            4'd8: result_0490 = (~((((b >> 2) | 14'd12176) - ((~14'd9142) - (b * 14'd9644))) ? (a ? ((b >> 1) ? (a ^ a) : 6171) : 3537) : 4809));
            
            4'd9: result_0490 = (((b + 14'd14505) - (14'd9778 * (14'd14516 & (b * a)))) + b);
            
            4'd10: result_0490 = (b >> 2);
            
            4'd11: result_0490 = (14'd1474 * (((14'd7565 * b) * ((a | b) * (14'd14736 | a))) - (((b ^ 14'd7499) ? (14'd11192 ? b : 5742) : 6844) ? ((~a) - (14'd1750 + 14'd15903)) : 4517)));
            
            default: result_0490 = 14'd10519;
        endcase
    end

endmodule
        