
module simple_alu_0818(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0818
);

    always @(*) begin
        case(op)
            
            4'd0: result_0818 = (b | a);
            
            4'd1: result_0818 = (((a | (~14'd6374)) - (((14'd7908 ^ a) << 3) ? (b + 14'd7376) : 7020)) * ((((14'd539 << 1) & 14'd15993) ? ((14'd6064 ^ 14'd1821) + (b - 14'd10414)) : 3508) >> 3));
            
            4'd2: result_0818 = ((b >> 2) - a);
            
            4'd3: result_0818 = (((((14'd3019 + b) >> 2) | (b - (a & 14'd2343))) * (((b << 2) | (a - 14'd7933)) & (~14'd10110))) ^ ((a >> 2) ^ (14'd4650 >> 1)));
            
            4'd4: result_0818 = ((a >> 1) & 14'd299);
            
            4'd5: result_0818 = ((14'd12084 | (14'd8321 - a)) * ((((14'd3306 - 14'd11269) * 14'd16344) | (14'd7082 - (b >> 1))) * 14'd2555));
            
            4'd6: result_0818 = (a ^ (14'd7895 >> 2));
            
            4'd7: result_0818 = ((14'd2733 + a) | 14'd7547);
            
            4'd8: result_0818 = (((((14'd3981 ? 14'd10455 : 748) | (14'd6827 ? a : 15480)) * ((14'd6288 & b) - (a * 14'd11092))) >> 2) * (a * (b * 14'd10015)));
            
            4'd9: result_0818 = (((b & ((14'd11021 ^ a) & 14'd181)) * a) + ((14'd9246 + 14'd350) | (14'd9892 + (14'd12846 & a))));
            
            4'd10: result_0818 = (a >> 1);
            
            4'd11: result_0818 = (a >> 3);
            
            4'd12: result_0818 = (((((14'd1437 >> 3) + (14'd11420 >> 1)) * (14'd4784 << 2)) >> 3) ? (14'd14782 ? ((14'd10279 | 14'd16342) & ((14'd6130 ? 14'd1015 : 12662) ^ a)) : 6112) : 11719);
            
            4'd13: result_0818 = (14'd11600 ? b : 6021);
            
            4'd14: result_0818 = (14'd15196 ^ ((((b >> 2) - (14'd7511 | b)) << 2) << 2));
            
            4'd15: result_0818 = ((~(~a)) ? 14'd3075 : 9342);
            
            default: result_0818 = 14'd13425;
        endcase
    end

endmodule
        