
module simple_alu_0327(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0327
);

    always @(*) begin
        case(op)
            
            4'd0: result_0327 = (14'd9437 | 14'd497);
            
            4'd1: result_0327 = (b + (~14'd9117));
            
            4'd2: result_0327 = ((b + (14'd14313 << 3)) >> 1);
            
            4'd3: result_0327 = ((14'd6794 + (((14'd9258 & 14'd8591) | (a - 14'd12647)) * b)) | ((~(14'd4835 * (~14'd11678))) << 3));
            
            4'd4: result_0327 = (~b);
            
            4'd5: result_0327 = ((~((~(14'd7464 ^ 14'd2434)) + ((14'd16204 + 14'd11452) ? (b >> 3) : 6219))) * ((b - 14'd5524) - (((14'd4596 ^ 14'd4733) - b) & (14'd13375 ^ (14'd10408 + a)))));
            
            4'd6: result_0327 = ((~(14'd3999 & ((14'd8398 | b) << 1))) & ((b & ((b * b) ^ (14'd6274 ^ a))) * (b - 14'd411)));
            
            4'd7: result_0327 = ((b - 14'd794) | 14'd10085);
            
            4'd8: result_0327 = (((((14'd11581 * 14'd3289) * (~14'd16337)) & 14'd15293) ? (14'd2806 << 1) : 6097) ? ((((14'd15480 + a) ? (14'd10114 ^ 14'd3926) : 14437) ? 14'd6126 : 866) ? b : 97) : 6192);
            
            4'd9: result_0327 = (14'd263 >> 1);
            
            4'd10: result_0327 = ((~14'd13686) ^ (((~14'd15751) | 14'd1400) ^ ((~(14'd6191 | a)) & ((a << 2) >> 3))));
            
            4'd11: result_0327 = (((((a >> 2) | 14'd8041) + (14'd1071 * (14'd6260 * 14'd9515))) - 14'd2898) >> 3);
            
            4'd12: result_0327 = (((((b ? 14'd11258 : 9922) | (14'd16340 & 14'd12925)) - 14'd2789) & (14'd2493 | (~14'd13562))) >> 3);
            
            4'd13: result_0327 = ((((a ? (a | a) : 3086) | 14'd10003) - (((b ? 14'd8112 : 7850) ^ (~b)) ^ 14'd6124)) | (14'd6770 >> 3));
            
            default: result_0327 = 14'd7814;
        endcase
    end

endmodule
        