
module simple_alu_0609(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0609
);

    always @(*) begin
        case(op)
            
            4'd0: result_0609 = ((~((b ? (14'd5216 ? 14'd300 : 15999) : 2856) ? b : 12492)) & (14'd9457 >> 2));
            
            4'd1: result_0609 = (14'd6731 - (~(((b >> 2) << 1) >> 1)));
            
            4'd2: result_0609 = ((~(14'd2392 << 1)) + (((14'd6049 + b) | ((~14'd10387) | b)) << 3));
            
            4'd3: result_0609 = (((((14'd7489 | a) & (14'd13824 ? 14'd3871 : 9491)) & 14'd3733) | ((b | (14'd5573 ? 14'd570 : 15582)) ? (14'd8447 ? 14'd6487 : 7243) : 11687)) - (((14'd7350 | (14'd12559 - 14'd14880)) - b) ^ (((~a) + 14'd3898) | (~(14'd14861 + 14'd8073)))));
            
            4'd4: result_0609 = ((((14'd13630 ^ (14'd6970 << 1)) | ((14'd13575 & b) << 1)) | (((14'd15168 ^ 14'd5660) + (a << 1)) >> 1)) & ((14'd12437 << 1) ^ (((a >> 1) ^ (14'd8152 >> 1)) | ((14'd2916 + 14'd2300) + (b ^ 14'd14168)))));
            
            4'd5: result_0609 = (((((a | 14'd15627) ^ (14'd14278 << 1)) << 2) ? (~(14'd11219 ^ (a & a))) : 3458) - 14'd933);
            
            4'd6: result_0609 = (14'd15980 ^ 14'd11896);
            
            4'd7: result_0609 = (((((14'd10041 << 3) * (14'd11387 - a)) >> 1) >> 1) - b);
            
            default: result_0609 = 14'd15421;
        endcase
    end

endmodule
        