
module simple_alu_0136(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0136
);

    always @(*) begin
        case(op)
            
            4'd0: result_0136 = (14'd2648 ? ((14'd12847 & 14'd11646) + (b ^ ((b ^ 14'd1921) ^ (14'd5111 ? 14'd8535 : 14291)))) : 16032);
            
            4'd1: result_0136 = (((~((~a) | (~14'd9535))) - (14'd8050 << 3)) >> 1);
            
            4'd2: result_0136 = (((((14'd5642 ^ a) | (14'd1141 << 3)) ? ((a << 3) + (14'd718 * 14'd4929)) : 13479) + ((14'd4120 ^ (14'd12975 - 14'd7338)) * ((14'd3644 >> 1) + a))) << 3);
            
            4'd3: result_0136 = (((14'd8717 | ((a * b) * (14'd1010 | 14'd7529))) ^ 14'd4556) ? ((((a - 14'd7542) | a) | (a >> 2)) ^ (((14'd14821 & 14'd10306) * (14'd1325 ^ 14'd13056)) | ((b >> 2) + (14'd6518 * b)))) : 4642);
            
            4'd4: result_0136 = ((b + 14'd6824) * (((14'd13662 & (b + b)) & 14'd13629) - (14'd8387 - ((14'd5289 & 14'd8696) ^ (b ^ 14'd4073)))));
            
            4'd5: result_0136 = ((b ? (((14'd1419 + a) ^ (a << 3)) ? (14'd9726 ^ 14'd9892) : 5675) : 9036) >> 2);
            
            4'd6: result_0136 = ((((~(14'd8644 & 14'd13106)) << 3) ? (((14'd6934 - 14'd15998) | (14'd8722 * b)) & (14'd12072 & (14'd12811 & 14'd6877))) : 9252) - ((~((~14'd14521) >> 3)) | 14'd2963));
            
            4'd7: result_0136 = ((((14'd8263 | (14'd288 >> 2)) | b) | ((a * 14'd13458) >> 2)) * ((~((14'd2953 ^ b) | (b ^ 14'd2433))) * ((14'd12537 ? 14'd1104 : 3128) * ((14'd6026 - a) ^ 14'd9321))));
            
            4'd8: result_0136 = (14'd7415 | (a ^ (((b - 14'd15972) - (14'd3109 & 14'd4783)) ? a : 4970)));
            
            4'd9: result_0136 = (14'd10494 | ((~(b & (a << 2))) ? (14'd6562 << 3) : 4605));
            
            4'd10: result_0136 = (((14'd10967 * ((a - 14'd6500) ? (a & 14'd6675) : 68)) - a) ? (a + b) : 7388);
            
            4'd11: result_0136 = (((((14'd11292 ^ 14'd5364) + b) << 3) | (((a | 14'd83) + (b * 14'd16218)) ? a : 11536)) ^ (~(14'd14657 & 14'd889)));
            
            default: result_0136 = a;
        endcase
    end

endmodule
        