
module simple_alu_0078(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0078
);

    always @(*) begin
        case(op)
            
            4'd0: result_0078 = (((((14'd13626 - 14'd3488) & (14'd5617 * 14'd13082)) + ((14'd6490 & 14'd8452) - (14'd6457 & 14'd2857))) << 2) + (((~(b | 14'd945)) >> 2) << 2));
            
            4'd1: result_0078 = (((14'd11701 * ((14'd13892 ? 14'd8397 : 5525) ? (14'd5145 ? 14'd9309 : 13454) : 14410)) | ((14'd16305 + (~14'd13716)) & ((14'd6991 * 14'd13206) & (14'd7151 + 14'd4453)))) & ((b & ((a | 14'd4108) - (b + 14'd15427))) ? (((a | a) - 14'd9928) & (14'd14751 * 14'd4964)) : 11060));
            
            4'd2: result_0078 = (((b << 2) ^ (((14'd14380 * a) ? 14'd7140 : 3210) << 3)) & ((((14'd1984 ? 14'd3789 : 8905) >> 1) - 14'd570) ^ 14'd3578));
            
            4'd3: result_0078 = (~(~((b >> 3) & ((a - a) << 3))));
            
            4'd4: result_0078 = (b | (14'd12739 & a));
            
            4'd5: result_0078 = ((14'd1060 & (((14'd8608 - 14'd11947) ? (a * 14'd15145) : 8214) | ((a ? b : 12806) >> 3))) * 14'd4968);
            
            4'd6: result_0078 = ((14'd7204 ^ (a + (14'd2426 ^ (a & 14'd6845)))) << 2);
            
            4'd7: result_0078 = (((((14'd5740 + a) << 2) & b) ? b : 10246) | ((~(14'd13187 + (14'd5804 << 3))) ? (14'd14309 ? 14'd4193 : 10912) : 12808));
            
            4'd8: result_0078 = (((((b ^ 14'd57) << 1) ^ (14'd9596 << 1)) & ((~(~14'd11125)) ^ (b | (14'd2405 * a)))) * 14'd10013);
            
            4'd9: result_0078 = (~14'd2097);
            
            4'd10: result_0078 = ((~((b ? 14'd3268 : 15509) & (~14'd9476))) << 1);
            
            default: result_0078 = 14'd14362;
        endcase
    end

endmodule
        