
module simple_alu_0619(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0619
);

    always @(*) begin
        case(op)
            
            4'd0: result_0619 = ((a * b) >> 3);
            
            4'd1: result_0619 = (b >> 3);
            
            4'd2: result_0619 = (((((a | 14'd4379) - 14'd12231) << 1) << 2) * ((((14'd4474 ? 14'd7152 : 10094) * (a ^ 14'd11770)) & (a + a)) ^ a));
            
            4'd3: result_0619 = (~(14'd1717 ^ (a & a)));
            
            4'd4: result_0619 = ((14'd14404 * (((14'd9589 - b) >> 1) - (14'd12593 | (~14'd14077)))) ? (b - ((~(14'd15147 | a)) << 2)) : 9495);
            
            4'd5: result_0619 = (((b >> 2) << 2) & 14'd1577);
            
            4'd6: result_0619 = ((14'd9467 << 2) ^ ((~((b * b) | b)) + 14'd4300));
            
            4'd7: result_0619 = (((14'd12157 ? ((a | b) - (~b)) : 10756) - (14'd7964 | ((b ^ b) - 14'd5762))) + (~(((~14'd3851) << 1) ? a : 416)));
            
            4'd8: result_0619 = ((((14'd7466 ^ (14'd7709 << 2)) << 3) | (14'd10857 >> 1)) ? (~14'd5648) : 6885);
            
            4'd9: result_0619 = ((14'd15851 & ((14'd9124 ? (b >> 3) : 13089) ^ ((14'd15991 << 2) << 2))) >> 3);
            
            4'd10: result_0619 = (((((14'd14847 >> 3) & (a * 14'd5289)) | (~(14'd966 << 3))) + ((~(14'd15609 - 14'd4673)) ^ ((14'd3006 & a) << 2))) >> 3);
            
            4'd11: result_0619 = (((14'd13314 >> 3) ^ (((14'd9274 * b) - (14'd6324 << 3)) ? (14'd13716 ? (b + 14'd3941) : 14076) : 6144)) * ((((14'd12675 | 14'd8226) ? a : 11915) * ((a | a) & (14'd9752 & b))) << 1));
            
            4'd12: result_0619 = (14'd14692 & b);
            
            4'd13: result_0619 = (((((14'd14535 ^ a) | (a | 14'd2134)) << 1) * (14'd5539 ? 14'd8979 : 15450)) >> 2);
            
            default: result_0619 = 14'd13518;
        endcase
    end

endmodule
        