
module simple_alu_0136(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0136
);

    always @(*) begin
        case(op)
            
            4'd0: result_0136 = ((((a - a) ? (12'd3322 << 2) : 1864) >> 2) + ((~(12'd3482 + b)) ^ (12'd3825 << 1)));
            
            4'd1: result_0136 = ((((b << 3) << 3) ? a : 1498) >> 3);
            
            4'd2: result_0136 = (12'd871 - (((12'd351 >> 2) - 12'd3634) ? (~(a & 12'd1861)) : 3043));
            
            4'd3: result_0136 = ((a ^ a) ? (((12'd2596 | 12'd2325) << 1) * (~b)) : 1431);
            
            4'd4: result_0136 = (((b - a) - ((b ^ 12'd3095) - (12'd2694 | 12'd3230))) & (~(b ? (a + 12'd3929) : 631)));
            
            4'd5: result_0136 = ((12'd1334 ? 12'd3643 : 3174) + (a * (a + (b * a))));
            
            4'd6: result_0136 = (~(a ^ (b | (12'd3061 << 3))));
            
            4'd7: result_0136 = (((~(a ? b : 232)) + ((b ^ a) ? 12'd1028 : 1537)) << 1);
            
            4'd8: result_0136 = (((~b) * ((~b) ^ (12'd3420 ^ b))) ^ (((b << 2) >> 1) & ((~b) << 3)));
            
            4'd9: result_0136 = (a ? ((12'd2601 << 1) ? 12'd1404 : 3610) : 2527);
            
            4'd10: result_0136 = (((b & 12'd748) * (a * 12'd2046)) << 2);
            
            4'd11: result_0136 = ((((~a) * (b + b)) | (b + (12'd3895 << 2))) << 1);
            
            4'd12: result_0136 = ((((12'd2653 >> 3) * (~12'd1966)) << 2) >> 1);
            
            default: result_0136 = 12'd3164;
        endcase
    end

endmodule
        