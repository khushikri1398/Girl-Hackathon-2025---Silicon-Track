
module simple_alu_0751(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0751
);

    always @(*) begin
        case(op)
            
            4'd0: result_0751 = (~(((a | 14'd12028) - (14'd8807 ? (14'd6410 & 14'd5175) : 13208)) | (14'd3683 - ((b * b) ? (a >> 1) : 16365))));
            
            4'd1: result_0751 = ((((~14'd8076) ^ ((14'd934 >> 3) << 2)) & (a ? b : 14426)) >> 3);
            
            4'd2: result_0751 = (14'd9017 << 3);
            
            4'd3: result_0751 = ((14'd9758 * (b ^ ((14'd6890 ? 14'd9263 : 13148) ? (~b) : 8470))) << 2);
            
            4'd4: result_0751 = ((b << 1) << 3);
            
            4'd5: result_0751 = ((14'd470 + (((b >> 2) * (b << 2)) << 3)) & (a * ((14'd10863 + 14'd5385) & 14'd16034)));
            
            4'd6: result_0751 = (((~b) ^ ((14'd251 << 2) << 2)) << 3);
            
            4'd7: result_0751 = (((((14'd1920 << 3) << 3) ^ 14'd3703) >> 1) | ((((14'd5618 >> 1) + (b & 14'd7578)) & ((b >> 3) ^ (a >> 1))) | b));
            
            4'd8: result_0751 = (((((a >> 3) * (14'd10294 ^ 14'd9074)) + (a << 1)) + (((14'd3205 << 3) >> 1) ^ 14'd6200)) >> 1);
            
            4'd9: result_0751 = ((~14'd9346) & ((((14'd14419 | 14'd119) >> 3) + 14'd4146) >> 1));
            
            4'd10: result_0751 = (14'd15380 | 14'd3920);
            
            4'd11: result_0751 = (((((14'd10549 << 2) ^ 14'd15953) ^ b) << 2) ^ (a << 1));
            
            default: result_0751 = b;
        endcase
    end

endmodule
        