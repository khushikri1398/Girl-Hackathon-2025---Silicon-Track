
module simple_alu_0120(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0120
);

    always @(*) begin
        case(op)
            
            4'd0: result_0120 = (~((((b & 14'd14838) + (14'd1632 << 1)) * ((14'd7936 + a) >> 3)) >> 1));
            
            4'd1: result_0120 = ((((14'd399 >> 3) << 1) + ((~(14'd15702 * 14'd3327)) << 1)) + ((14'd9217 * ((14'd11096 * 14'd799) ? (14'd7351 - 14'd7139) : 13612)) >> 2));
            
            4'd2: result_0120 = ((((14'd2824 - (14'd5603 << 3)) >> 2) | (((b * 14'd3097) - a) << 2)) - b);
            
            4'd3: result_0120 = (~a);
            
            4'd4: result_0120 = (~14'd2016);
            
            4'd5: result_0120 = (((((14'd8696 + b) | 14'd3419) << 3) - (14'd3358 + ((14'd13733 - a) ^ (~b)))) ^ ((~(14'd12175 ^ b)) * 14'd6896));
            
            4'd6: result_0120 = (14'd13940 ^ (((b >> 1) ^ ((14'd5614 - b) - (14'd2329 ? 14'd3970 : 1838))) & ((14'd6171 << 1) << 2)));
            
            4'd7: result_0120 = (((14'd2881 | ((14'd16278 >> 2) | 14'd5874)) ? 14'd14506 : 15672) & 14'd4100);
            
            4'd8: result_0120 = (~14'd5208);
            
            4'd9: result_0120 = (~(14'd12918 ^ ((14'd8690 << 2) ? 14'd3234 : 3294)));
            
            4'd10: result_0120 = (((((~b) * (14'd4358 - a)) - ((14'd2874 << 2) * (14'd13299 - a))) << 2) + ((((~a) | b) | (14'd6198 >> 3)) >> 1));
            
            4'd11: result_0120 = (((((14'd14324 * 14'd5237) << 2) ? a : 11600) + (~((a << 1) - (14'd10791 >> 1)))) >> 1);
            
            4'd12: result_0120 = (((b ? (~(a & a)) : 2597) | (((~b) ? (b & 14'd2403) : 2124) >> 2)) | (((b << 3) * ((14'd8696 ^ 14'd3083) ? (14'd14967 | 14'd2462) : 1377)) * (~((14'd5644 ^ 14'd3238) ^ (14'd11673 | a)))));
            
            4'd13: result_0120 = ((14'd9084 * ((14'd5477 | a) ? (~(14'd12574 + 14'd1570)) : 4210)) | (b | ((14'd4627 | 14'd11080) >> 3)));
            
            4'd14: result_0120 = ((b | (~b)) * (b >> 2));
            
            4'd15: result_0120 = (((14'd9657 | a) ? a : 9484) ^ (~((~(14'd6009 | 14'd7922)) ^ 14'd5124)));
            
            default: result_0120 = a;
        endcase
    end

endmodule
        