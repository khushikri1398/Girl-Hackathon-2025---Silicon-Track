
module simple_alu_0370(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0370
);

    always @(*) begin
        case(op)
            
            4'd0: result_0370 = (((a ^ ((a & 14'd12330) - (14'd3450 - 14'd1563))) >> 2) >> 1);
            
            4'd1: result_0370 = (((((b ^ 14'd2205) ? (a >> 1) : 3987) + ((a * 14'd8792) ^ (14'd4483 + 14'd658))) & 14'd10607) - ((((14'd14355 | a) << 3) ^ 14'd6721) & ((~(14'd8971 ? b : 11094)) >> 3)));
            
            4'd2: result_0370 = ((~(~((~14'd9513) & 14'd7806))) << 3);
            
            4'd3: result_0370 = ((~((a | 14'd3431) - ((14'd10486 ^ a) - (14'd7198 ^ 14'd10504)))) + (((~(~14'd13198)) + 14'd15604) + b));
            
            4'd4: result_0370 = (~(14'd12072 - ((b << 2) - 14'd4959)));
            
            4'd5: result_0370 = (((14'd3067 >> 2) + (b - (~(a ^ 14'd1354)))) * 14'd7539);
            
            4'd6: result_0370 = (14'd10439 ? (((b + (14'd10561 >> 2)) | (a + 14'd6491)) + ((14'd1914 - (14'd15027 >> 2)) + ((14'd5354 * 14'd63) >> 1))) : 5961);
            
            4'd7: result_0370 = (((((b & b) << 1) & ((a - b) + (b - 14'd1100))) - (((14'd7035 ? 14'd3171 : 10873) ^ (14'd2111 ^ 14'd15621)) * ((~14'd8612) * 14'd3990))) & 14'd8541);
            
            4'd8: result_0370 = ((((a >> 3) | 14'd7332) + (14'd4044 + ((14'd5771 ? 14'd8050 : 4988) & (14'd15963 >> 2)))) ^ (((a & (~a)) | (b ^ b)) >> 3));
            
            4'd9: result_0370 = ((a + (14'd16088 | 14'd5469)) - a);
            
            4'd10: result_0370 = (((((14'd9717 * 14'd9884) - (a + 14'd9434)) >> 2) | (((14'd2324 + b) * (a >> 2)) - ((14'd11317 - a) | (b >> 1)))) << 2);
            
            4'd11: result_0370 = (((((14'd2389 & 14'd15003) + (~14'd3386)) + (~14'd12130)) * (14'd8367 ? (14'd11027 ? (~a) : 13641) : 8597)) - ((((a ? a : 11373) ^ (b * 14'd7242)) ? ((14'd4369 >> 2) & (14'd16074 + a)) : 14702) | (14'd10497 + 14'd10787)));
            
            default: result_0370 = 14'd15018;
        endcase
    end

endmodule
        