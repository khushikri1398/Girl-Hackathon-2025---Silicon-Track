
module simple_alu_0486(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0486
);

    always @(*) begin
        case(op)
            
            4'd0: result_0486 = (a - ((((~b) ^ (14'd10074 + a)) << 2) * (((a * b) >> 3) * ((b & a) >> 3))));
            
            4'd1: result_0486 = (((((14'd15188 ^ 14'd12550) & (14'd6170 & b)) ^ 14'd5594) >> 3) + ((b << 1) & 14'd3691));
            
            4'd2: result_0486 = ((14'd9103 << 2) | ((((14'd6125 & b) ? (~a) : 11533) >> 3) << 3));
            
            4'd3: result_0486 = (b * a);
            
            4'd4: result_0486 = ((14'd4016 + (((14'd9700 + a) ? (b + 14'd786) : 2047) ? ((a >> 3) & (~a)) : 255)) >> 2);
            
            4'd5: result_0486 = (~(((14'd51 ? (14'd13477 ? a : 12191) : 240) * 14'd9665) & (((a << 2) + (b << 2)) >> 1)));
            
            4'd6: result_0486 = ((((~(a | 14'd11254)) ^ 14'd263) ? ((14'd13275 ^ (~14'd2463)) ? ((b * 14'd5240) ^ (14'd11245 >> 2)) : 7692) : 5990) << 1);
            
            4'd7: result_0486 = ((14'd15843 - (a & (~(~14'd3399)))) & (((14'd2838 + (14'd651 + b)) | 14'd228) >> 3));
            
            4'd8: result_0486 = ((14'd5401 | (((b << 1) & b) * ((14'd8969 ? 14'd12988 : 10318) >> 3))) | (14'd14471 ^ (((14'd16204 ^ b) ^ (14'd15103 ^ 14'd4025)) ? 14'd15394 : 15752)));
            
            4'd9: result_0486 = ((((~(~14'd13933)) * ((~14'd7630) & b)) | ((~(14'd6041 << 3)) - 14'd4749)) + a);
            
            4'd10: result_0486 = ((b << 3) ^ (14'd14571 >> 3));
            
            4'd11: result_0486 = (14'd11525 & ((((14'd1952 ? 14'd14631 : 4174) - (~a)) >> 2) | (b << 2)));
            
            default: result_0486 = 14'd12288;
        endcase
    end

endmodule
        