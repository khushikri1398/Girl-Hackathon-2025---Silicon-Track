
module simple_alu_0620(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0620
);

    always @(*) begin
        case(op)
            
            4'd0: result_0620 = (((b | ((14'd4519 ? b : 15810) ? (b & b) : 9486)) * (((14'd8583 + 14'd15492) & (b * 14'd12612)) * 14'd1977)) - a);
            
            4'd1: result_0620 = ((b * (14'd10152 << 1)) - ((((14'd4234 >> 2) + (~14'd11886)) + ((a * 14'd3402) >> 3)) + a));
            
            4'd2: result_0620 = ((14'd10219 - ((a ? (b ? 14'd5800 : 522) : 5026) << 3)) - (~(14'd8196 | a)));
            
            4'd3: result_0620 = ((((b - 14'd11974) ? ((14'd11101 << 3) | (~14'd6005)) : 8590) << 1) & ((b + (14'd11797 ^ (a & a))) - 14'd10451));
            
            4'd4: result_0620 = ((14'd15088 + (((a | 14'd16048) >> 2) + ((14'd5596 * b) ? (14'd6095 | b) : 12220))) | 14'd6517);
            
            4'd5: result_0620 = (14'd14739 >> 2);
            
            4'd6: result_0620 = (((a << 2) ^ (((14'd8784 + 14'd8054) ^ (14'd13753 * 14'd3443)) - ((14'd13035 * 14'd9399) ? (~14'd7041) : 15526))) << 1);
            
            4'd7: result_0620 = (14'd5818 - (~(((b ? 14'd2370 : 1316) >> 2) | ((14'd13583 << 2) | (14'd15449 & b)))));
            
            4'd8: result_0620 = ((b >> 3) ^ ((b ? ((b ^ 14'd5094) + a) : 2461) ^ (((a & 14'd2783) ^ (a & a)) * (14'd14082 & (a - b)))));
            
            4'd9: result_0620 = (((((14'd3016 ^ 14'd13738) | (b | a)) << 3) ^ (((a ? a : 6003) * (14'd11908 ^ 14'd14297)) + ((14'd16114 * 14'd5760) << 3))) | ((((a ? 14'd10863 : 8646) ^ b) * a) - a));
            
            4'd10: result_0620 = ((((b - (a - 14'd702)) * ((b - a) * (b ^ 14'd11501))) - (14'd14804 ? ((~b) >> 2) : 920)) ^ 14'd11783);
            
            4'd11: result_0620 = ((~((14'd4542 + 14'd2823) & ((14'd12954 - 14'd13200) - (14'd16063 >> 1)))) << 1);
            
            4'd12: result_0620 = (((14'd10617 >> 2) - (~((~14'd15827) ? (14'd15588 << 3) : 7409))) & b);
            
            4'd13: result_0620 = (((((~a) * 14'd4402) & ((14'd4164 * 14'd3875) | (a << 1))) & b) << 2);
            
            default: result_0620 = b;
        endcase
    end

endmodule
        