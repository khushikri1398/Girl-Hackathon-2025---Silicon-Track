
module simple_alu_0103(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0103
);

    always @(*) begin
        case(op)
            
            4'd0: result_0103 = (((((14'd519 << 1) | b) & ((14'd4754 * 14'd2098) | 14'd3726)) & (((14'd7735 * b) ^ 14'd7548) * (~(14'd11520 ? a : 8113)))) - 14'd6145);
            
            4'd1: result_0103 = (14'd16060 >> 1);
            
            4'd2: result_0103 = (((((14'd14675 - 14'd9220) * (14'd571 - 14'd15096)) ^ b) & 14'd1751) + (a | a));
            
            4'd3: result_0103 = (((b | ((b & 14'd10563) << 2)) & (14'd2992 - 14'd10647)) - ((((14'd6889 ? 14'd13354 : 2763) >> 1) << 2) - (((a + 14'd3478) - (14'd6353 - 14'd8801)) ^ 14'd5793)));
            
            4'd4: result_0103 = (~((((14'd15039 ? 14'd7149 : 12438) - (14'd14818 & 14'd14131)) | 14'd14404) + ((14'd4112 - (a | 14'd9928)) + 14'd1050)));
            
            4'd5: result_0103 = (~14'd5289);
            
            4'd6: result_0103 = (14'd4956 >> 3);
            
            4'd7: result_0103 = (a * (((~(b ? 14'd15278 : 5967)) >> 2) ^ 14'd15800));
            
            4'd8: result_0103 = (((~(14'd3802 + (b * 14'd9311))) ? (((a & a) ^ (14'd7548 + a)) << 1) : 5310) + ((14'd12019 | ((14'd11728 * 14'd5608) * (14'd8429 | 14'd5843))) >> 1));
            
            default: result_0103 = b;
        endcase
    end

endmodule
        