
module simple_alu_0303(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0303
);

    always @(*) begin
        case(op)
            
            4'd0: result_0303 = (a ^ (14'd1960 & a));
            
            4'd1: result_0303 = (14'd2877 * (b - ((~(14'd1602 ^ b)) ? ((b << 2) << 3) : 15209)));
            
            4'd2: result_0303 = ((~14'd4924) * (((14'd6373 ^ (14'd6520 - 14'd9551)) & 14'd15632) >> 2));
            
            4'd3: result_0303 = (14'd8341 << 2);
            
            4'd4: result_0303 = (((a & 14'd15354) ? (((14'd14133 - 14'd3720) - 14'd10174) + 14'd11607) : 8287) & 14'd3781);
            
            4'd5: result_0303 = (14'd13354 ^ (a >> 2));
            
            4'd6: result_0303 = (((14'd13529 >> 1) >> 1) & b);
            
            4'd7: result_0303 = (14'd7172 << 2);
            
            4'd8: result_0303 = (14'd10892 >> 2);
            
            4'd9: result_0303 = ((14'd2539 + 14'd15226) | 14'd16229);
            
            4'd10: result_0303 = ((b | ((14'd4124 << 1) >> 3)) << 1);
            
            4'd11: result_0303 = ((b & ((14'd1397 - (14'd13033 | 14'd5219)) + ((b | 14'd12423) ? (~14'd4702) : 14268))) << 3);
            
            4'd12: result_0303 = (14'd11453 << 3);
            
            default: result_0303 = b;
        endcase
    end

endmodule
        