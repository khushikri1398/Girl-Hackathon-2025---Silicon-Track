
module simple_alu_0294(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0294
);

    always @(*) begin
        case(op)
            
            4'd0: result_0294 = (~(14'd7840 - ((a << 3) ^ ((a ? a : 7954) ? (b ^ 14'd15842) : 12427))));
            
            4'd1: result_0294 = (((((b | a) ^ (b | a)) ? 14'd13346 : 56) + ((~14'd14932) ^ ((14'd11014 - 14'd324) ? (a & b) : 3417))) * ((14'd7080 ^ ((14'd8729 ? 14'd13510 : 10076) & a)) & (((a * 14'd5415) ^ (b | 14'd8774)) * (a + (14'd8995 << 2)))));
            
            4'd2: result_0294 = (((14'd14843 ^ ((14'd7283 << 2) >> 3)) ? 14'd3855 : 164) >> 3);
            
            4'd3: result_0294 = (((((b - 14'd2346) & 14'd3156) ? b : 5862) * (a ? ((b & 14'd1505) << 3) : 10118)) & (((14'd8755 | 14'd13471) - ((14'd7889 + 14'd6497) & (~14'd884))) << 1));
            
            4'd4: result_0294 = (((14'd7031 - ((a ^ 14'd15019) | (14'd15853 ^ a))) ^ (((b << 1) << 1) & 14'd2094)) ? 14'd8774 : 11014);
            
            4'd5: result_0294 = ((14'd4289 ^ b) ^ ((b ^ 14'd6718) >> 1));
            
            4'd6: result_0294 = (((14'd9642 << 3) - b) ? 14'd2956 : 14929);
            
            default: result_0294 = b;
        endcase
    end

endmodule
        