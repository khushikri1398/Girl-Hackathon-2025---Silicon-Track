
module simple_alu_0584(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0584
);

    always @(*) begin
        case(op)
            
            4'd0: result_0584 = ((((14'd3855 << 2) >> 1) ^ (~(14'd2913 | 14'd5060))) | ((((14'd14695 << 3) & (14'd3014 >> 3)) ^ (14'd3830 & 14'd14490)) - (~((14'd12313 * 14'd2143) & (b | a)))));
            
            4'd1: result_0584 = (14'd1979 ? (a << 1) : 1491);
            
            4'd2: result_0584 = ((14'd15027 - b) - ((~b) & 14'd16109));
            
            4'd3: result_0584 = (b >> 2);
            
            4'd4: result_0584 = (14'd618 - (((b >> 2) + 14'd3368) * 14'd7867));
            
            4'd5: result_0584 = (a ? 14'd2744 : 13557);
            
            4'd6: result_0584 = ((b | ((b * (14'd9654 & 14'd8564)) << 1)) << 2);
            
            4'd7: result_0584 = (a & (14'd825 ^ b));
            
            4'd8: result_0584 = ((14'd2500 - (~((14'd13310 << 1) - (14'd2893 + b)))) | ((14'd15225 | 14'd486) | (((a - 14'd11088) ^ 14'd1916) + ((14'd15682 | b) + (14'd3939 >> 3)))));
            
            4'd9: result_0584 = (((((14'd7290 ? 14'd13691 : 15010) - (14'd3275 - 14'd3446)) & 14'd14002) & (((14'd6731 >> 3) >> 3) ^ ((14'd10254 << 3) ^ (14'd4763 << 3)))) ^ (14'd1071 ? a : 8377));
            
            4'd10: result_0584 = ((14'd3410 & (~(~(a << 3)))) ? (14'd4055 + 14'd3649) : 7927);
            
            4'd11: result_0584 = (((((14'd1312 - b) ^ 14'd11008) | (a - (14'd9604 >> 1))) << 1) - 14'd14997);
            
            4'd12: result_0584 = ((((~14'd11860) * ((14'd10999 >> 3) >> 1)) >> 2) - (a ? (14'd4119 * ((~b) ^ (14'd6861 - 14'd12707))) : 710));
            
            4'd13: result_0584 = (14'd7555 * b);
            
            4'd14: result_0584 = (((b * ((14'd1476 << 1) | (14'd8485 & 14'd749))) ^ (((14'd1591 | 14'd9566) >> 3) * ((14'd12349 ^ b) | (b + 14'd16046)))) >> 3);
            
            default: result_0584 = 14'd722;
        endcase
    end

endmodule
        