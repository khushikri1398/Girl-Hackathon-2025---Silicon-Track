
module simple_alu_0082(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0082
);

    always @(*) begin
        case(op)
            
            4'd0: result_0082 = (b >> 2);
            
            4'd1: result_0082 = (~(14'd3876 << 2));
            
            4'd2: result_0082 = (14'd13543 | (14'd11685 - a));
            
            4'd3: result_0082 = (((b >> 3) + ((~(14'd5135 << 1)) >> 1)) | ((((a & b) & (14'd5246 | 14'd7839)) * ((14'd5618 & 14'd3238) ^ (a >> 3))) + 14'd14622));
            
            4'd4: result_0082 = (14'd10346 & (((b | (14'd782 - 14'd7049)) ^ (b - (~b))) | b));
            
            4'd5: result_0082 = (((((14'd12882 - a) ^ 14'd3224) << 1) & 14'd11465) ? 14'd9194 : 11632);
            
            4'd6: result_0082 = (b - 14'd14971);
            
            4'd7: result_0082 = (~((((14'd7511 - 14'd9583) ? (14'd15163 ^ b) : 8259) >> 2) * 14'd11719));
            
            4'd8: result_0082 = ((((~(a * 14'd13051)) & ((14'd15126 + 14'd11387) * 14'd9620)) * ((a & (14'd13370 >> 1)) | 14'd7514)) - a);
            
            4'd9: result_0082 = (b - (~(a | a)));
            
            4'd10: result_0082 = ((a + (~14'd4245)) >> 3);
            
            4'd11: result_0082 = ((b & 14'd15184) | ((14'd13323 << 1) | (14'd11936 - ((14'd927 + a) | (~a)))));
            
            4'd12: result_0082 = (((14'd12625 | (b ^ (14'd5325 + 14'd10748))) + (~(14'd13629 - a))) - ((b * (a >> 2)) | b));
            
            4'd13: result_0082 = (14'd15612 ? 14'd12192 : 11881);
            
            default: result_0082 = 14'd363;
        endcase
    end

endmodule
        