
module simple_alu_0395(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0395
);

    always @(*) begin
        case(op)
            
            4'd0: result_0395 = ((a * (~((14'd1824 << 1) << 3))) ^ (a ? a : 8685));
            
            4'd1: result_0395 = ((((b ^ 14'd7444) - (~(~14'd6301))) << 3) - (b ? (((a + 14'd13484) + 14'd15948) ^ ((14'd4158 >> 2) * b)) : 4519));
            
            4'd2: result_0395 = (14'd4511 ^ (((~(b >> 2)) << 1) ? (((14'd15111 & 14'd12429) - (a & 14'd11955)) & b) : 4727));
            
            4'd3: result_0395 = (((((b ? 14'd5987 : 3386) ^ 14'd13396) * ((14'd6025 + a) << 3)) - 14'd8194) ? ((((14'd12223 | 14'd3817) >> 1) << 2) ^ (~((14'd9037 << 1) + b))) : 11329);
            
            4'd4: result_0395 = (14'd15835 ^ (~((14'd4554 ? (b & 14'd2336) : 5694) ^ (~(14'd12340 << 2)))));
            
            default: result_0395 = 14'd4536;
        endcase
    end

endmodule
        