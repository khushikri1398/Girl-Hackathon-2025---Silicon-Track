
module simple_alu_0491(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0491
);

    always @(*) begin
        case(op)
            
            4'd0: result_0491 = (14'd11683 ? b : 10022);
            
            4'd1: result_0491 = (a * b);
            
            4'd2: result_0491 = ((((a ? (14'd494 * 14'd14844) : 726) ? ((14'd8745 ? 14'd13475 : 5864) ? 14'd433 : 11453) : 14672) - (((14'd3078 | b) ? (14'd8285 << 2) : 15956) + (~(14'd3980 ? b : 12143)))) - (((a - (a * a)) - 14'd15468) & (14'd12294 | 14'd14435)));
            
            4'd3: result_0491 = ((~(((14'd15651 << 1) ^ (14'd16263 - 14'd13276)) * (14'd10130 * (14'd4557 ? 14'd12343 : 1392)))) | (~((14'd11072 + (a | 14'd11175)) << 2)));
            
            4'd4: result_0491 = ((14'd15448 & (14'd8514 * a)) >> 3);
            
            4'd5: result_0491 = (((14'd3047 * b) + 14'd7188) * (14'd4375 | b));
            
            4'd6: result_0491 = ((14'd7887 - (~(14'd11122 ^ (14'd744 - 14'd5666)))) << 1);
            
            4'd7: result_0491 = (((((a * b) >> 2) | ((14'd4736 >> 1) << 2)) + (((14'd7318 & 14'd9487) & (14'd10827 << 1)) | (~14'd13269))) * ((14'd3490 + (~(14'd9927 << 1))) & 14'd329));
            
            4'd8: result_0491 = ((b & 14'd337) | (~((a + (14'd15555 * b)) ? ((14'd11553 ^ 14'd12591) ^ (14'd7482 + a)) : 1391)));
            
            4'd9: result_0491 = (a ? b : 10579);
            
            4'd10: result_0491 = (b ^ ((((b - a) ? (~a) : 8090) - 14'd3421) | (b ? (~14'd7170) : 1772)));
            
            4'd11: result_0491 = (((~14'd9997) & (((a << 1) + (a & 14'd3610)) ^ ((a - b) << 1))) << 1);
            
            4'd12: result_0491 = (b + (~(a | ((b - 14'd10934) + (14'd1443 * a)))));
            
            4'd13: result_0491 = ((14'd7324 + (a | 14'd8658)) ? (~14'd6863) : 1736);
            
            4'd14: result_0491 = (14'd4266 * ((((~b) << 3) - (14'd5387 - (14'd330 + a))) >> 3));
            
            default: result_0491 = b;
        endcase
    end

endmodule
        