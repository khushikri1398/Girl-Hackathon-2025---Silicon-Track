
module simple_alu_0300(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0300
);

    always @(*) begin
        case(op)
            
            4'd0: result_0300 = ((((12'd4037 ? 12'd279 : 2438) >> 2) | ((~12'd1656) & 12'd3373)) ^ 12'd3140);
            
            4'd1: result_0300 = ((((~b) >> 3) * ((12'd541 ? a : 3728) & 12'd3981)) >> 3);
            
            4'd2: result_0300 = (12'd502 | 12'd1579);
            
            4'd3: result_0300 = ((((a >> 1) + b) ? 12'd1526 : 1205) - 12'd2390);
            
            4'd4: result_0300 = ((((12'd1478 + 12'd2243) + (12'd4045 << 1)) + ((a >> 3) ^ (12'd1461 * a))) | 12'd3375);
            
            4'd5: result_0300 = ((((12'd3223 * a) * (12'd840 * 12'd2684)) & b) >> 2);
            
            4'd6: result_0300 = ((((12'd3050 ^ 12'd2669) >> 3) & ((12'd3121 | 12'd1789) ? (a * 12'd1621) : 588)) >> 3);
            
            4'd7: result_0300 = ((((12'd2464 ? 12'd375 : 884) ^ (12'd2653 ^ 12'd3373)) | 12'd3630) & 12'd3225);
            
            4'd8: result_0300 = ((~a) | (((12'd963 + 12'd2651) - (b * 12'd3151)) ^ ((12'd298 - 12'd2017) - (12'd4048 + a))));
            
            4'd9: result_0300 = ((((12'd2963 >> 2) ^ (b ^ 12'd3537)) & (12'd80 * b)) & 12'd217);
            
            4'd10: result_0300 = (~(((12'd1297 >> 3) << 1) + (12'd822 | (12'd3110 | 12'd739))));
            
            4'd11: result_0300 = (((~(a | 12'd3993)) | ((b ? a : 2468) ? (~b) : 3714)) | (((a & 12'd1977) ^ 12'd2078) ^ (12'd863 << 2)));
            
            4'd12: result_0300 = (((12'd2249 | (b ? b : 608)) * 12'd2887) ^ 12'd3512);
            
            default: result_0300 = 12'd769;
        endcase
    end

endmodule
        