
module simple_alu_0051(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0051
);

    always @(*) begin
        case(op)
            
            4'd0: result_0051 = (14'd12132 ^ ((14'd15601 * ((b >> 2) >> 3)) | ((b + b) + b)));
            
            4'd1: result_0051 = (((((~14'd10360) >> 3) + ((14'd7619 >> 1) * 14'd5123)) >> 3) | a);
            
            4'd2: result_0051 = (((((b ^ b) | (b ? 14'd4459 : 9776)) & ((a - 14'd442) | (a * a))) >> 2) & ((((b & a) * (14'd13856 >> 2)) | ((a & 14'd2666) ^ 14'd3041)) + (((a + b) ? 14'd7907 : 11366) + ((14'd3414 >> 1) ^ (14'd13224 - 14'd3331)))));
            
            4'd3: result_0051 = (b ^ (((14'd1444 ^ (a | 14'd6587)) ? ((b - 14'd13016) | b) : 4099) * (((a + a) - 14'd9049) + ((a ? b : 14953) ? 14'd14878 : 11851))));
            
            4'd4: result_0051 = ((b - (a + 14'd1184)) + ((~(a - (b ? b : 4875))) | (14'd13974 | a)));
            
            4'd5: result_0051 = ((14'd6905 << 3) * 14'd6295);
            
            4'd6: result_0051 = (b * ((((14'd16017 + a) << 3) << 2) ^ (b ^ a)));
            
            4'd7: result_0051 = (((b ^ (14'd13519 ? (a ? a : 13046) : 12646)) << 2) + a);
            
            default: result_0051 = 14'd2280;
        endcase
    end

endmodule
        