
module simple_alu_0381(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0381
);

    always @(*) begin
        case(op)
            
            4'd0: result_0381 = (((((b ^ b) << 2) + ((14'd1717 * b) + (a + b))) & (((14'd1760 ? 14'd9588 : 230) & (a | 14'd14691)) * (14'd15657 & (b << 2)))) ^ (((a << 1) ^ ((14'd818 & 14'd14934) * (a * a))) * b));
            
            4'd1: result_0381 = (((((a - 14'd15661) - a) ? ((a | 14'd16251) | (14'd15390 ^ b)) : 3257) & 14'd9221) ? ((14'd3383 ? a : 15976) ? 14'd14436 : 14492) : 16381);
            
            4'd2: result_0381 = (b >> 3);
            
            4'd3: result_0381 = (((~b) * (((b ? 14'd935 : 1374) ^ (a & 14'd224)) + ((14'd7379 - 14'd12900) + (14'd808 - b)))) & ((((b ^ 14'd10169) & (b & 14'd8869)) - ((a | a) - 14'd5745)) & (((a << 2) ? a : 13841) >> 1)));
            
            4'd4: result_0381 = (((((14'd1723 * b) * 14'd11533) & (a - (b << 2))) | (((14'd15011 + 14'd5936) << 2) >> 1)) - (~a));
            
            4'd5: result_0381 = (((((b << 3) * 14'd8278) << 3) ^ (b >> 2)) | (((a >> 1) | (14'd8864 >> 2)) * 14'd2096));
            
            4'd6: result_0381 = (((((b - 14'd13089) & (14'd5180 >> 2)) << 2) ^ b) | (a * (14'd6882 << 1)));
            
            4'd7: result_0381 = (14'd16376 >> 1);
            
            default: result_0381 = 14'd4633;
        endcase
    end

endmodule
        