
module simple_alu_0177(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0177
);

    always @(*) begin
        case(op)
            
            4'd0: result_0177 = ((14'd10333 ^ 14'd15276) * ((14'd14679 ^ ((~a) ^ (~14'd15626))) >> 3));
            
            4'd1: result_0177 = (~(14'd3779 - (((14'd4161 ? 14'd9337 : 971) << 2) - a)));
            
            4'd2: result_0177 = (b - (((b + 14'd14028) << 3) & (~(b - 14'd4906))));
            
            4'd3: result_0177 = (((~((14'd10129 ^ b) & (b << 2))) >> 3) * b);
            
            4'd4: result_0177 = (14'd3322 >> 3);
            
            4'd5: result_0177 = (a + (14'd9833 ? (((14'd5283 & a) | 14'd1411) * 14'd10723) : 12262));
            
            4'd6: result_0177 = ((b << 3) << 2);
            
            4'd7: result_0177 = (~(14'd9098 | (((14'd8218 ? 14'd15462 : 1494) ^ 14'd12924) ? 14'd14580 : 9580)));
            
            4'd8: result_0177 = ((((14'd2749 - 14'd4825) + ((14'd6110 | b) ^ 14'd2552)) * (((a >> 1) ? 14'd11715 : 1382) & b)) | (b + (((b ? 14'd5689 : 2383) << 3) ? ((a ? b : 6069) - (14'd15026 ? 14'd9804 : 16220)) : 12277)));
            
            4'd9: result_0177 = (((b & a) >> 2) >> 3);
            
            4'd10: result_0177 = ((14'd4462 + (14'd4514 & ((14'd7739 << 2) - b))) & (~a));
            
            4'd11: result_0177 = (14'd6010 & 14'd3377);
            
            4'd12: result_0177 = ((14'd2043 << 1) * (14'd468 & ((~(14'd5092 >> 3)) - (~(a & 14'd553)))));
            
            4'd13: result_0177 = (((((b | a) + (14'd12625 * a)) * ((14'd3740 + 14'd10301) ? b : 15650)) >> 3) >> 3);
            
            4'd14: result_0177 = ((((~(14'd16381 + a)) * (14'd4942 >> 1)) | 14'd5358) + (~14'd5712));
            
            default: result_0177 = 14'd6186;
        endcase
    end

endmodule
        