
module simple_alu_0363(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0363
);

    always @(*) begin
        case(op)
            
            4'd0: result_0363 = ((~a) + 14'd9518);
            
            4'd1: result_0363 = (((14'd2051 ? ((14'd9404 << 1) ? (14'd2804 ? 14'd13905 : 14476) : 16201) : 12252) * (((a ^ 14'd11924) >> 2) - ((a - 14'd4546) >> 2))) | 14'd525);
            
            4'd2: result_0363 = ((~(((14'd9281 ? a : 3409) << 3) - (14'd9237 * (14'd739 >> 2)))) * (14'd3276 >> 1));
            
            4'd3: result_0363 = (((14'd6914 - ((a | 14'd5900) ^ (14'd15471 >> 1))) ? a : 6214) >> 3);
            
            4'd4: result_0363 = ((((~a) - ((a & 14'd13635) | (a & 14'd16250))) ^ 14'd1032) + (a >> 2));
            
            4'd5: result_0363 = (a & 14'd11313);
            
            4'd6: result_0363 = (((14'd11533 & b) * 14'd11704) * ((((14'd4880 ^ 14'd9627) & a) & 14'd992) >> 3));
            
            4'd7: result_0363 = ((((14'd11993 + (a * b)) - (a ? (a + a) : 5946)) << 1) >> 3);
            
            4'd8: result_0363 = (~(b >> 3));
            
            default: result_0363 = 14'd13399;
        endcase
    end

endmodule
        