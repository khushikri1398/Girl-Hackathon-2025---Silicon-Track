
module simple_alu_0497(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0497
);

    always @(*) begin
        case(op)
            
            4'd0: result_0497 = ((b ? (~((~14'd13470) - (14'd1152 * 14'd9986))) : 13782) | ((~((14'd10925 << 2) - (a | 14'd12449))) >> 1));
            
            4'd1: result_0497 = (~((b >> 2) ^ (~(14'd9540 ^ (14'd3759 >> 2)))));
            
            4'd2: result_0497 = ((14'd12194 ^ ((a ^ (14'd5625 + b)) - (14'd11722 ? (b ^ 14'd9575) : 8436))) ^ b);
            
            4'd3: result_0497 = (((~((14'd5561 | a) - b)) & (b & ((a >> 3) & 14'd15773))) | 14'd9636);
            
            4'd4: result_0497 = ((((~(b | b)) | ((14'd11925 + 14'd4517) >> 2)) + 14'd10914) << 1);
            
            4'd5: result_0497 = ((14'd5504 + (((b ^ b) - (b * a)) ^ 14'd456)) + (b + (((14'd8197 ? 14'd9422 : 5085) ? (b & 14'd4498) : 11353) - ((14'd14985 ? 14'd4807 : 8112) - (a | 14'd3372)))));
            
            4'd6: result_0497 = ((((a | (b * 14'd2713)) ? ((14'd11168 + a) - (14'd6880 * 14'd8008)) : 16141) ^ (14'd13139 + ((14'd15900 - a) + (a << 1)))) | (((14'd1046 & (~14'd5875)) * (~14'd15806)) << 1));
            
            4'd7: result_0497 = ((~(~((14'd6866 - 14'd6651) ? (a >> 2) : 9925))) | ((14'd10508 >> 3) * 14'd2960));
            
            default: result_0497 = a;
        endcase
    end

endmodule
        