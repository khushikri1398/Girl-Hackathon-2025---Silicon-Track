
module simple_alu_0272(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0272
);

    always @(*) begin
        case(op)
            
            4'd0: result_0272 = (a - ((14'd1002 | ((14'd12933 * 14'd8089) ? (14'd14278 >> 2) : 8467)) ? (((14'd5697 << 3) - (14'd3350 << 3)) * ((14'd11393 ? a : 10974) | (14'd6193 - b))) : 13329));
            
            4'd1: result_0272 = ((((14'd879 + (14'd12973 | 14'd10238)) | ((14'd4367 + 14'd11842) ^ (14'd8023 & a))) ? (((14'd8395 | b) >> 2) << 2) : 13786) ^ (((14'd8434 << 3) - ((a << 3) << 2)) << 2));
            
            4'd2: result_0272 = (14'd6871 * ((((14'd8425 - 14'd7591) & (a & 14'd9540)) ^ ((b ^ b) ? 14'd16297 : 5194)) + ((~(~b)) ? ((b | 14'd13633) >> 3) : 1144)));
            
            4'd3: result_0272 = (((((b + a) >> 3) * ((~14'd8972) | (14'd13703 >> 3))) ? (14'd3081 - (a ? b : 11087)) : 10397) << 3);
            
            4'd4: result_0272 = (((((14'd2190 * 14'd9970) + (14'd12107 ? a : 15435)) - ((b >> 3) + a)) - a) ^ b);
            
            4'd5: result_0272 = (((((b >> 1) >> 2) ^ ((b ? a : 2452) | (14'd6374 * 14'd4082))) ? ((14'd3966 << 2) ? (b - a) : 6224) : 12090) << 3);
            
            4'd6: result_0272 = (~((((a ^ a) << 2) >> 3) - ((~14'd6818) & 14'd10164)));
            
            4'd7: result_0272 = ((14'd13163 + (a + ((a * b) * (14'd13173 & b)))) | ((14'd8847 << 3) >> 2));
            
            4'd8: result_0272 = ((~(14'd15820 ^ ((a - 14'd16224) | (14'd10964 >> 1)))) ^ ((((b - 14'd12196) + 14'd3504) + b) ^ (((b & 14'd586) >> 2) ^ b)));
            
            default: result_0272 = b;
        endcase
    end

endmodule
        