
module simple_alu_0245(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0245
);

    always @(*) begin
        case(op)
            
            4'd0: result_0245 = ((~14'd3057) & a);
            
            4'd1: result_0245 = ((~14'd11257) >> 1);
            
            4'd2: result_0245 = (((((14'd1642 ? 14'd11436 : 6182) - (~14'd5149)) ? ((a ^ a) << 2) : 12995) * 14'd12480) - (b - (((14'd3149 ^ b) + a) << 3)));
            
            4'd3: result_0245 = (((~14'd14550) >> 3) * b);
            
            4'd4: result_0245 = (14'd6552 & ((b * (14'd1280 - (a | 14'd14648))) ^ (~(14'd9274 - a))));
            
            4'd5: result_0245 = (b | ((((14'd4965 ? 14'd2227 : 8203) | (14'd881 - 14'd6883)) - ((b * 14'd15227) & (b & b))) | ((14'd10120 >> 1) * ((14'd6085 & a) & (b << 2)))));
            
            4'd6: result_0245 = (((~(~a)) | (((a + 14'd5482) + (14'd11215 >> 3)) ? (b ^ 14'd2770) : 10855)) ? (14'd9211 << 3) : 7563);
            
            4'd7: result_0245 = (((((a ? b : 7772) - (14'd6998 * a)) - (~14'd10286)) & b) | 14'd7626);
            
            4'd8: result_0245 = ((~((~14'd9096) & ((14'd6522 ? 14'd8721 : 2629) ^ (~14'd15178)))) ? ((((14'd4159 - 14'd9809) | (b - 14'd9846)) + ((14'd15649 << 3) - (a - 14'd4509))) >> 2) : 242);
            
            4'd9: result_0245 = (((((a ^ 14'd11792) ? (a ^ a) : 8534) << 1) - (((14'd12358 | 14'd6415) ? (a ? 14'd4993 : 1798) : 15032) * (14'd11900 - (a >> 1)))) - (a * (14'd12813 | (~14'd7804))));
            
            4'd10: result_0245 = (~(b | (((b ^ a) & a) >> 1)));
            
            4'd11: result_0245 = (~(((14'd6696 | (14'd6960 - 14'd12149)) >> 1) - 14'd5777));
            
            4'd12: result_0245 = (14'd11747 << 2);
            
            4'd13: result_0245 = (14'd13267 & ((~((14'd4481 & a) << 3)) & 14'd4789));
            
            default: result_0245 = 14'd16022;
        endcase
    end

endmodule
        