
module simple_alu_0803(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0803
);

    always @(*) begin
        case(op)
            
            4'd0: result_0803 = (14'd2019 >> 3);
            
            4'd1: result_0803 = (((14'd13031 & 14'd14247) | (14'd11098 << 2)) * ((((14'd2534 ^ 14'd15186) ^ (14'd6889 & 14'd5325)) + 14'd3909) | (((14'd14983 + a) + (14'd13646 >> 1)) << 2)));
            
            4'd2: result_0803 = (((((14'd3289 - b) ? (b ? 14'd3711 : 1877) : 3060) - 14'd8476) + (~((14'd4056 ^ 14'd7138) * (14'd8441 * a)))) << 2);
            
            4'd3: result_0803 = (((14'd3713 ? (14'd788 << 1) : 12763) & (((14'd1383 * 14'd15736) * (14'd15014 >> 1)) * (~b))) ? 14'd15876 : 4340);
            
            4'd4: result_0803 = (14'd5347 ? 14'd2540 : 2899);
            
            4'd5: result_0803 = (14'd11657 + (14'd10076 >> 1));
            
            4'd6: result_0803 = (14'd9649 ? 14'd5658 : 16363);
            
            4'd7: result_0803 = (14'd16144 ^ ((((14'd609 + b) & (a & a)) ^ ((14'd4349 ^ 14'd16308) ? (14'd9404 ? 14'd13840 : 4892) : 10394)) >> 1));
            
            4'd8: result_0803 = ((14'd3420 | a) ? (14'd6669 | (((14'd7396 + a) * 14'd6224) ^ 14'd8862)) : 5442);
            
            4'd9: result_0803 = ((14'd13802 - 14'd4051) ? (((14'd12602 + (14'd13143 | 14'd4244)) ? ((a + 14'd414) | 14'd10379) : 8773) | 14'd12155) : 6223);
            
            4'd10: result_0803 = (((((a >> 3) * (a ? a : 325)) - b) * (b | ((14'd6499 & b) * (~14'd9978)))) - ((a ^ ((a * b) | (a >> 1))) * (14'd13556 + (b >> 2))));
            
            4'd11: result_0803 = (((((14'd11877 ^ 14'd294) >> 1) - a) - b) << 2);
            
            4'd12: result_0803 = (((((14'd6195 ? 14'd5441 : 1427) >> 2) ? ((a ^ 14'd15978) + (a ? 14'd15351 : 2078)) : 3303) ^ b) | b);
            
            default: result_0803 = a;
        endcase
    end

endmodule
        