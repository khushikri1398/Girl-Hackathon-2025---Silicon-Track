
module simple_alu_0905(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0905
);

    always @(*) begin
        case(op)
            
            4'd0: result_0905 = ((((14'd13307 << 3) - b) ? (((14'd9101 - 14'd6863) >> 1) ? ((b + b) ? (14'd12002 ? 14'd5166 : 10859) : 2981) : 16293) : 12757) | (~((14'd7345 | (a - a)) ? (~(14'd15321 - b)) : 11467)));
            
            4'd1: result_0905 = (14'd534 & 14'd15011);
            
            4'd2: result_0905 = (((((~a) << 2) ^ a) ? (b ? a : 695) : 10275) >> 1);
            
            4'd3: result_0905 = (14'd11769 ^ ((a & 14'd1330) + ((~(b | 14'd6571)) | (14'd15137 << 1))));
            
            4'd4: result_0905 = (a & ((((b | 14'd9697) - 14'd4892) << 2) & (((~b) & 14'd1767) - ((~14'd9556) + (b ^ a)))));
            
            4'd5: result_0905 = (((((14'd7982 + 14'd15942) ^ (14'd3027 >> 2)) & 14'd695) ^ 14'd228) + 14'd3931);
            
            4'd6: result_0905 = (~14'd10418);
            
            4'd7: result_0905 = (((~((a - a) - (b * 14'd14499))) | (~((14'd6810 >> 3) ^ (~14'd3119)))) + (a ? 14'd5956 : 7331));
            
            4'd8: result_0905 = (14'd9260 + (~(14'd6569 << 1)));
            
            4'd9: result_0905 = (14'd6713 - ((~14'd8539) | (14'd10218 - (a | (14'd5201 ^ 14'd1380)))));
            
            4'd10: result_0905 = (((14'd13793 - 14'd11027) >> 2) >> 3);
            
            default: result_0905 = 14'd4550;
        endcase
    end

endmodule
        