
module simple_alu_0745(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0745
);

    always @(*) begin
        case(op)
            
            4'd0: result_0745 = ((((b & 14'd1694) ? ((a >> 1) + (b - b)) : 15637) * (((14'd4048 - 14'd13393) ^ (14'd14201 ? 14'd9509 : 7919)) ? ((14'd2203 ? 14'd7387 : 15056) >> 3) : 434)) + 14'd9079);
            
            4'd1: result_0745 = (((((a & a) | a) + 14'd7455) & (((14'd14737 & 14'd4590) | (a | a)) * 14'd8185)) + a);
            
            4'd2: result_0745 = ((((b >> 1) ? ((b - 14'd8946) - (14'd6496 ^ 14'd8264)) : 10046) + (14'd13588 >> 2)) ? (14'd190 - (((a ^ 14'd3210) ^ (~b)) + ((b << 3) ^ 14'd3862))) : 10932);
            
            4'd3: result_0745 = (((((a & 14'd15940) | (14'd5091 ^ 14'd13807)) ? (b * a) : 3248) << 2) + a);
            
            4'd4: result_0745 = (b & (((b - (14'd279 | b)) - 14'd14958) & (~((a ? b : 10692) ? (14'd11923 << 3) : 10284))));
            
            4'd5: result_0745 = (((((14'd6530 * 14'd14579) >> 1) + a) * (((14'd7007 ? b : 7414) * (a >> 1)) - (14'd575 ? (14'd8309 << 2) : 13072))) | 14'd3968);
            
            4'd6: result_0745 = ((14'd13431 << 3) ^ 14'd10050);
            
            4'd7: result_0745 = (14'd10258 ^ (~a));
            
            4'd8: result_0745 = (a ? (14'd7299 >> 2) : 7453);
            
            4'd9: result_0745 = ((14'd3662 & (14'd14547 ? ((a ? a : 11242) << 2) : 2004)) - ((((14'd12326 ? b : 13056) - a) >> 2) + ((14'd13028 ? (b ^ b) : 6699) >> 1)));
            
            4'd10: result_0745 = (((b >> 2) << 1) & (~14'd5422));
            
            4'd11: result_0745 = (14'd11834 >> 2);
            
            4'd12: result_0745 = ((~(~((b & 14'd4449) ^ (14'd5013 - 14'd5731)))) >> 3);
            
            4'd13: result_0745 = (a << 3);
            
            default: result_0745 = a;
        endcase
    end

endmodule
        