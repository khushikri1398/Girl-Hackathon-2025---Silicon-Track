
module simple_alu_0296(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0296
);

    always @(*) begin
        case(op)
            
            4'd0: result_0296 = ((a >> 2) * ((((14'd7528 << 3) ^ 14'd3142) | ((a << 3) | (a * a))) & (b + ((14'd9658 >> 3) | (14'd600 | 14'd8705)))));
            
            4'd1: result_0296 = (14'd328 & a);
            
            4'd2: result_0296 = (14'd8545 ^ ((~((b * 14'd13893) ? (~b) : 5526)) << 2));
            
            4'd3: result_0296 = ((a ^ (((14'd1271 << 3) ^ (14'd2880 << 2)) ? a : 717)) + ((((14'd13367 ^ 14'd1964) >> 3) - b) >> 2));
            
            4'd4: result_0296 = ((14'd3147 - (((14'd1389 << 1) & 14'd297) ? (14'd15528 | (b - 14'd16091)) : 10757)) ? ((((~14'd6598) << 2) >> 2) | ((~a) << 2)) : 3927);
            
            4'd5: result_0296 = (14'd7935 | ((((~b) << 3) + 14'd12152) * (((14'd8658 | 14'd145) ^ (~14'd12416)) >> 3)));
            
            4'd6: result_0296 = (((((b | 14'd9387) * (14'd3609 >> 1)) ^ 14'd13336) & (((14'd4199 | a) - 14'd3859) >> 1)) | 14'd4078);
            
            4'd7: result_0296 = (b & 14'd13447);
            
            4'd8: result_0296 = (~14'd14437);
            
            4'd9: result_0296 = (((14'd15858 - ((b & 14'd4700) ? (b + 14'd7016) : 2472)) >> 3) * 14'd1304);
            
            default: result_0296 = 14'd10796;
        endcase
    end

endmodule
        