
module simple_alu_0636(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0636
);

    always @(*) begin
        case(op)
            
            4'd0: result_0636 = (((b * ((~14'd10000) ? (b - 14'd11413) : 11573)) >> 3) * a);
            
            4'd1: result_0636 = (((14'd11109 << 1) ^ (((14'd9563 & 14'd14548) ^ b) ? ((14'd145 | a) | (14'd1693 - 14'd7993)) : 1352)) << 1);
            
            4'd2: result_0636 = ((b & a) << 1);
            
            4'd3: result_0636 = ((~((a >> 3) - ((14'd16269 ^ 14'd15160) >> 3))) ? (14'd6642 * (~((a << 3) * (a & 14'd1876)))) : 2016);
            
            4'd4: result_0636 = (~((((14'd10156 | 14'd13876) ? (14'd11294 + b) : 11533) + ((b | 14'd10831) ? (14'd3398 + 14'd4693) : 8502)) * 14'd1827));
            
            4'd5: result_0636 = (~((((b * 14'd3123) - (a * 14'd5043)) + b) + (((14'd13304 * 14'd15070) << 2) ? ((a | b) & 14'd8378) : 15969)));
            
            4'd6: result_0636 = ((b & 14'd10570) + (b + ((14'd15120 + (b & b)) * ((~14'd4021) & (14'd2447 * a)))));
            
            4'd7: result_0636 = ((14'd6044 ^ ((~(~14'd14065)) + ((14'd4448 - b) ^ (a | 14'd10903)))) ? 14'd4136 : 14736);
            
            4'd8: result_0636 = (((14'd15278 << 1) - 14'd5198) & 14'd12534);
            
            4'd9: result_0636 = (((14'd12751 | ((14'd1056 | 14'd12500) & (~14'd3604))) >> 2) & 14'd10085);
            
            4'd10: result_0636 = (14'd15681 | (14'd11657 + b));
            
            4'd11: result_0636 = (((~(14'd6015 & b)) >> 1) - ((((14'd14893 | 14'd8827) - (b * b)) >> 3) | ((14'd1193 ? (14'd11593 & 14'd3395) : 12684) ? ((14'd12104 ^ a) & (b + a)) : 5161)));
            
            4'd12: result_0636 = (((a ^ 14'd299) ? (((14'd13664 ? 14'd11325 : 5472) >> 3) | ((b ^ 14'd13805) * (14'd9341 | 14'd13442))) : 7325) & b);
            
            4'd13: result_0636 = ((((b >> 1) << 3) * (((a >> 1) * b) & (14'd3485 >> 1))) >> 3);
            
            4'd14: result_0636 = (((~((14'd14186 + 14'd2945) << 3)) + 14'd8640) - (((14'd13459 | (14'd11468 - a)) * ((14'd14179 | b) & (14'd14858 ^ b))) - (14'd1411 & (~14'd15695))));
            
            4'd15: result_0636 = (14'd4242 ^ 14'd5161);
            
            default: result_0636 = 14'd7688;
        endcase
    end

endmodule
        