
module simple_alu_0098(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0098
);

    always @(*) begin
        case(op)
            
            4'd0: result_0098 = (b ^ ((((a << 2) << 1) & (b ^ b)) ^ b));
            
            4'd1: result_0098 = ((14'd14312 ? a : 3533) ? (14'd10492 >> 3) : 9936);
            
            4'd2: result_0098 = (((((b ^ a) + 14'd2958) * (14'd5359 >> 2)) & (~((14'd13530 >> 2) | (14'd7026 & b)))) * ((a >> 3) ? 14'd15426 : 6952));
            
            4'd3: result_0098 = (((~((~14'd14250) & b)) >> 1) * (((~(a | a)) ? 14'd9338 : 7977) + (((14'd7663 - 14'd3271) * (14'd12009 + 14'd13552)) + (b & a))));
            
            4'd4: result_0098 = (14'd2374 & (14'd5078 * 14'd6937));
            
            4'd5: result_0098 = ((((~(a ? 14'd5943 : 3340)) & ((14'd14680 ? b : 15140) ^ 14'd11118)) + 14'd8936) * (b * (((b + 14'd13966) + (~14'd9817)) ? (~(a + 14'd12815)) : 4705)));
            
            4'd6: result_0098 = (((~((14'd14372 ^ b) << 1)) ? 14'd2735 : 8489) * (b - (((14'd10187 - 14'd7864) >> 3) >> 3)));
            
            4'd7: result_0098 = ((~(((14'd5810 & 14'd9795) & (14'd10862 | 14'd15375)) | (~(a - a)))) + 14'd6055);
            
            4'd8: result_0098 = (((a & (a - 14'd15777)) + 14'd7404) ? ((14'd11573 - ((14'd6435 * 14'd8893) ^ a)) ^ (14'd8732 | (~(14'd101 ^ 14'd5253)))) : 12599);
            
            4'd9: result_0098 = ((((b ? (14'd2979 - 14'd9753) : 8263) | (b ? (14'd14794 & 14'd15594) : 15972)) << 2) >> 1);
            
            default: result_0098 = 14'd65;
        endcase
    end

endmodule
        