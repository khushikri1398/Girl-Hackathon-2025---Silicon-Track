
module simple_alu_0866(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0866
);

    always @(*) begin
        case(op)
            
            4'd0: result_0866 = (((((14'd2842 << 3) & b) >> 3) & 14'd4526) ? a : 9776);
            
            4'd1: result_0866 = ((((14'd7777 & a) & 14'd15198) - (((~b) * (14'd8542 + 14'd13680)) ^ (~14'd11163))) ? ((((a ^ 14'd13550) ? a : 11749) - b) - (((14'd11475 & 14'd16268) ^ 14'd7581) * ((~b) - 14'd7453))) : 3770);
            
            4'd2: result_0866 = (((~(~(14'd14179 * 14'd15305))) >> 3) ? (((14'd9469 ^ (14'd6596 ? b : 12144)) << 2) >> 2) : 10035);
            
            4'd3: result_0866 = (b >> 2);
            
            4'd4: result_0866 = (((((a + 14'd377) | (14'd9417 * 14'd8594)) >> 2) + (~((14'd7747 & 14'd7581) | 14'd9060))) ^ ((14'd9282 + ((b ^ a) & (~a))) * (14'd8384 ^ b)));
            
            4'd5: result_0866 = (((14'd1509 << 1) ^ ((14'd4152 ^ (14'd1173 | b)) & ((a ? a : 15124) + (14'd8312 << 2)))) << 2);
            
            4'd6: result_0866 = (((14'd12451 + 14'd1755) >> 3) ^ (((14'd10573 << 1) & (~a)) + b));
            
            4'd7: result_0866 = (((((14'd4650 - a) + b) >> 2) ? (~a) : 9446) | (((14'd2860 << 1) ^ ((a ? a : 647) >> 1)) ^ a));
            
            4'd8: result_0866 = (~14'd857);
            
            4'd9: result_0866 = (~14'd8647);
            
            default: result_0866 = a;
        endcase
    end

endmodule
        