
module simple_alu_0314(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0314
);

    always @(*) begin
        case(op)
            
            4'd0: result_0314 = (((a + (~(14'd3535 ? 14'd3783 : 8834))) + (a - (~(b + a)))) * 14'd7538);
            
            4'd1: result_0314 = ((~((b << 1) & a)) * (14'd4338 * ((14'd16002 & (14'd7077 ? a : 8449)) & ((~14'd5770) & (a ? b : 3260)))));
            
            4'd2: result_0314 = (a * ((((a & 14'd8662) * (14'd4020 ? a : 11990)) << 1) | 14'd963));
            
            4'd3: result_0314 = ((~(14'd7515 ? b : 863)) ^ ((((b | 14'd3586) * (14'd14868 ? 14'd6039 : 6412)) * ((~14'd15403) ? (b | 14'd15809) : 7514)) + 14'd11372));
            
            4'd4: result_0314 = ((((14'd7556 | a) << 1) ? (((14'd5144 >> 2) + (14'd16337 | 14'd783)) & ((14'd12494 - b) ? 14'd3218 : 9035)) : 10310) >> 2);
            
            4'd5: result_0314 = ((14'd12420 >> 1) ^ (((14'd109 | (14'd673 + 14'd7372)) | (~(b * 14'd9202))) * (((14'd11375 >> 2) - (b * 14'd1645)) * ((14'd14636 >> 3) >> 2))));
            
            4'd6: result_0314 = (~(~((14'd12180 | 14'd10211) ^ (14'd15392 >> 2))));
            
            default: result_0314 = 14'd2539;
        endcase
    end

endmodule
        