
module simple_alu_0655(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0655
);

    always @(*) begin
        case(op)
            
            4'd0: result_0655 = (((14'd512 << 3) & (((14'd13062 ^ a) | (14'd8639 << 2)) ? ((14'd12690 >> 2) - (14'd14541 | a)) : 4307)) * 14'd6760);
            
            4'd1: result_0655 = ((a << 1) ? (~(((a & b) + (14'd7243 * a)) ? (~(14'd3535 & 14'd12041)) : 15725)) : 8361);
            
            4'd2: result_0655 = (((((14'd15756 ^ 14'd14350) << 3) << 3) + (((14'd5050 * b) ^ (a + 14'd9544)) << 1)) ? b : 11201);
            
            4'd3: result_0655 = ((b ^ (((a + b) << 3) ^ 14'd5389)) * ((14'd14116 - ((a - a) | (14'd9580 + 14'd884))) ? a : 10446));
            
            4'd4: result_0655 = (14'd2495 - b);
            
            4'd5: result_0655 = (14'd1642 * ((((14'd11313 & a) - (14'd8931 ^ a)) | ((14'd3119 - 14'd14207) << 3)) & (~(~(14'd12341 ? 14'd4849 : 10426)))));
            
            4'd6: result_0655 = (~14'd15794);
            
            4'd7: result_0655 = (((a << 3) << 1) & 14'd12984);
            
            4'd8: result_0655 = (~(14'd13697 & (((14'd11864 | 14'd7474) - (b >> 2)) ? ((14'd12637 + a) | (14'd8580 ? b : 12989)) : 11961)));
            
            4'd9: result_0655 = (14'd13511 + b);
            
            4'd10: result_0655 = (14'd9845 >> 2);
            
            4'd11: result_0655 = (14'd2856 & ((((~14'd480) * 14'd175) - ((a >> 2) >> 2)) + (~14'd11949)));
            
            4'd12: result_0655 = (14'd1199 << 2);
            
            default: result_0655 = 14'd8440;
        endcase
    end

endmodule
        