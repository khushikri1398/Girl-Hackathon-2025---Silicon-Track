
module simple_alu_0483(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0483
);

    always @(*) begin
        case(op)
            
            4'd0: result_0483 = ((((b + (14'd6006 | a)) & 14'd11544) | (((14'd620 ^ a) & (a >> 3)) >> 3)) - ((a ? ((a - 14'd4639) ? b : 16169) : 10566) ? (((14'd8637 | a) << 2) * ((14'd14303 & b) * (~14'd5024))) : 14754));
            
            4'd1: result_0483 = ((((~a) << 3) - (((~b) + (b & 14'd8309)) ^ ((b - 14'd1309) * (b * b)))) | (((~(b & 14'd12196)) >> 3) << 2));
            
            4'd2: result_0483 = ((((~(14'd4837 & 14'd9047)) >> 3) & ((~(~14'd1587)) + ((14'd3347 * a) << 2))) - ((14'd12880 + (a ^ b)) ? (((a ? 14'd12028 : 250) >> 1) * ((b ? a : 5431) ? (14'd999 * b) : 6458)) : 14087));
            
            4'd3: result_0483 = ((((~(14'd9475 * 14'd16287)) - ((a * 14'd11649) << 1)) ^ ((~(b + 14'd9743)) ? ((14'd10018 & a) ? (14'd6594 + 14'd6536) : 7411) : 2337)) ? ((((14'd11905 >> 2) & (a + 14'd9085)) * ((~b) ^ (14'd851 ? 14'd16344 : 5444))) >> 3) : 12137);
            
            4'd4: result_0483 = (~14'd11039);
            
            4'd5: result_0483 = (a * ((a ^ ((14'd7924 | 14'd1019) * (14'd4727 | 14'd11083))) * (14'd4682 >> 3)));
            
            4'd6: result_0483 = ((((14'd6704 | 14'd12918) ? b : 3637) ? 14'd10644 : 15529) & ((b << 3) - (b | ((b * b) * (14'd9439 << 1)))));
            
            default: result_0483 = b;
        endcase
    end

endmodule
        