
module simple_alu_0368(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0368
);

    always @(*) begin
        case(op)
            
            4'd0: result_0368 = (~(~(b + (b << 2))));
            
            4'd1: result_0368 = (~((((~14'd12619) >> 2) >> 1) & ((~(a - 14'd4152)) + (a << 1))));
            
            4'd2: result_0368 = (((((14'd7251 | b) ^ (14'd13198 << 3)) << 3) * 14'd7137) & ((((b | b) >> 1) ^ ((~14'd14742) ? (b | 14'd2085) : 10184)) - ((b & (14'd8173 << 3)) >> 2)));
            
            4'd3: result_0368 = (~(((~(14'd11783 | b)) >> 1) << 2));
            
            4'd4: result_0368 = (((((14'd10657 ^ 14'd2056) + 14'd9731) & 14'd2206) + (((14'd4408 ? 14'd14815 : 9621) >> 2) + (14'd5603 & 14'd11655))) ^ b);
            
            4'd5: result_0368 = (14'd4950 & (14'd11903 >> 3));
            
            4'd6: result_0368 = (14'd13694 + (b * ((~14'd16342) + ((b << 1) ^ (14'd10492 ^ 14'd3002)))));
            
            4'd7: result_0368 = ((a & 14'd15741) << 1);
            
            4'd8: result_0368 = ((14'd5419 * (14'd12479 ^ ((a ^ a) + 14'd10626))) & ((14'd6044 ? ((14'd5680 << 1) * 14'd5718) : 6660) << 3));
            
            4'd9: result_0368 = (14'd10977 ^ ((14'd377 - 14'd2428) & (b + (~(14'd8225 | 14'd15064)))));
            
            4'd10: result_0368 = ((14'd11168 | (((14'd13391 - 14'd15243) * (14'd9881 | 14'd15239)) | b)) << 2);
            
            4'd11: result_0368 = (((b + ((14'd15642 | 14'd3236) ^ (a >> 1))) >> 3) - 14'd15847);
            
            4'd12: result_0368 = (((((b >> 1) - (b - 14'd10551)) | (14'd15256 + (b ? b : 1031))) ^ 14'd12351) >> 1);
            
            4'd13: result_0368 = (((((~14'd724) >> 3) & (a + (14'd3476 - 14'd7184))) | ((14'd8997 << 3) * (~(14'd9429 | 14'd15173)))) - 14'd9041);
            
            default: result_0368 = 14'd12184;
        endcase
    end

endmodule
        