
module simple_alu_0561(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0561
);

    always @(*) begin
        case(op)
            
            4'd0: result_0561 = (((((~a) ^ 14'd16139) - ((14'd8733 - 14'd4685) + (a ^ a))) - (b & 14'd5724)) & ((14'd752 & ((b ^ 14'd14507) * 14'd11128)) | ((14'd12332 & (14'd168 ? 14'd7567 : 6799)) << 1)));
            
            4'd1: result_0561 = (((14'd1862 >> 1) ^ ((14'd14937 | 14'd7396) + ((a ? 14'd2294 : 6828) << 2))) & (b >> 2));
            
            4'd2: result_0561 = ((14'd8949 & ((~(14'd1898 ^ b)) | (14'd10052 | (a + 14'd5031)))) << 1);
            
            4'd3: result_0561 = (b - (~(14'd13927 | (a & (14'd8066 | b)))));
            
            4'd4: result_0561 = (((a << 1) * (((14'd14453 | 14'd5434) * (a ? 14'd11861 : 13680)) ? b : 15078)) - 14'd9106);
            
            4'd5: result_0561 = ((~(14'd10403 << 3)) ? ((((b ^ 14'd9655) * a) >> 1) ^ (14'd8267 | ((14'd15590 ? b : 781) << 3))) : 13064);
            
            4'd6: result_0561 = (~b);
            
            4'd7: result_0561 = (14'd8778 - ((14'd13178 & 14'd3507) << 1));
            
            4'd8: result_0561 = (((((~14'd2812) * 14'd6372) + a) ^ (((14'd13111 - 14'd6896) >> 2) * (~a))) ? (14'd15175 + (((14'd2206 ? a : 8677) - 14'd11737) & ((a - b) & b))) : 14429);
            
            4'd9: result_0561 = (((14'd1895 & ((b * 14'd4429) & (14'd11920 - 14'd7872))) + (b | ((14'd1312 >> 1) + 14'd13687))) ? ((((a ? 14'd7223 : 13648) * (a + 14'd2335)) ^ ((14'd14634 * 14'd11154) >> 2)) + 14'd813) : 13574);
            
            4'd10: result_0561 = (((((14'd2046 & 14'd2762) * (14'd5748 + b)) | ((a << 1) << 2)) + 14'd9839) | ((((a & 14'd3607) ^ (~a)) ? ((14'd10636 - b) + (14'd12677 | b)) : 13127) | (((14'd15828 ^ a) ? (14'd10295 + a) : 6453) & ((a | 14'd2557) & 14'd4060))));
            
            4'd11: result_0561 = ((a + b) >> 3);
            
            default: result_0561 = 14'd9341;
        endcase
    end

endmodule
        