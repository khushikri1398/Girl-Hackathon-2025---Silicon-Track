
module simple_alu_0656(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0656
);

    always @(*) begin
        case(op)
            
            4'd0: result_0656 = ((b | b) | 14'd1740);
            
            4'd1: result_0656 = ((((~(14'd5988 << 1)) - (a - a)) + (((14'd12566 | b) | a) * (b >> 1))) + (~(((14'd8805 | 14'd16066) | b) * ((a & a) | (b | 14'd12062)))));
            
            4'd2: result_0656 = (((a >> 1) << 1) >> 2);
            
            4'd3: result_0656 = ((~((a & b) - (14'd11425 | 14'd1844))) ^ ((b << 1) * (((a ? 14'd4515 : 13680) << 1) + ((14'd11128 >> 2) ? (14'd16364 * 14'd4350) : 13814))));
            
            4'd4: result_0656 = (~(14'd12456 | (~a)));
            
            4'd5: result_0656 = (((((b & 14'd9698) * 14'd865) & (14'd6685 ^ (14'd15195 | 14'd14353))) << 1) - ((((b & b) | 14'd5334) & ((14'd4226 - 14'd5609) << 3)) & 14'd11336));
            
            4'd6: result_0656 = ((~(((a ^ 14'd2016) + (14'd10131 << 2)) ^ 14'd16333)) - ((((b ? 14'd14997 : 5149) - 14'd12105) - 14'd8476) - (14'd5614 * ((a - 14'd10838) ? a : 472))));
            
            4'd7: result_0656 = (a & b);
            
            4'd8: result_0656 = (14'd10328 + (14'd11959 ^ 14'd13692));
            
            4'd9: result_0656 = (((a >> 2) | (~14'd10211)) * ((((~b) ^ (14'd8685 ^ b)) - a) & 14'd3874));
            
            default: result_0656 = a;
        endcase
    end

endmodule
        