
module simple_alu_0368(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0368
);

    always @(*) begin
        case(op)
            
            4'd0: result_0368 = (~((((a & 14'd12238) + 14'd8069) >> 1) >> 3));
            
            4'd1: result_0368 = (((14'd12774 & (14'd3495 + (b >> 1))) - b) & (~(~((14'd8591 - 14'd11464) & 14'd8872))));
            
            4'd2: result_0368 = (~14'd5750);
            
            4'd3: result_0368 = ((((14'd4395 << 3) * ((14'd6406 * 14'd463) | a)) + ((14'd14997 >> 3) << 2)) << 2);
            
            4'd4: result_0368 = (~((a & a) ? (((14'd16065 * b) * (14'd9357 ^ 14'd10130)) | (~(14'd872 ^ b))) : 9055));
            
            4'd5: result_0368 = (14'd7103 | 14'd4083);
            
            4'd6: result_0368 = (~((((a | a) * (~b)) * ((14'd10366 ^ 14'd13233) + 14'd13293)) << 3));
            
            4'd7: result_0368 = (((b - b) - b) | 14'd9810);
            
            4'd8: result_0368 = (~(((~(b + 14'd6016)) << 2) | b));
            
            4'd9: result_0368 = (((~((a ^ 14'd5762) ^ 14'd14251)) + (14'd15018 | (14'd5130 << 1))) >> 1);
            
            4'd10: result_0368 = (~(14'd1310 - (((14'd14614 ^ a) + (14'd8101 + 14'd8585)) ^ ((a | 14'd11423) + a))));
            
            4'd11: result_0368 = (14'd3520 * (b << 2));
            
            4'd12: result_0368 = (14'd14553 * ((((b - 14'd14853) ^ (14'd16018 & 14'd15604)) >> 1) ? ((~(a ^ 14'd9071)) | (~14'd13308)) : 4943));
            
            default: result_0368 = b;
        endcase
    end

endmodule
        