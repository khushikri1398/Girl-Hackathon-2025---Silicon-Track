
module simple_alu_0337(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0337
);

    always @(*) begin
        case(op)
            
            4'd0: result_0337 = ((14'd2858 * (b | a)) & (b * (((a - 14'd122) ? (14'd3999 >> 1) : 6697) | ((14'd7484 & 14'd13649) - (~b)))));
            
            4'd1: result_0337 = (14'd8682 ^ ((~14'd1100) << 3));
            
            4'd2: result_0337 = ((~(14'd9022 ^ ((a + b) * (14'd1758 ^ a)))) - ((~14'd13071) ^ (((14'd8469 ^ 14'd13795) | (~14'd2050)) >> 3)));
            
            4'd3: result_0337 = (((((~b) + (a << 2)) | 14'd2766) + 14'd3505) - ((((14'd14500 & 14'd15610) * (14'd10841 + 14'd10451)) & (a << 3)) ? 14'd12224 : 4398));
            
            4'd4: result_0337 = (((((14'd4055 >> 1) | 14'd7380) >> 3) ^ 14'd469) - ((a & a) ? ((~(14'd7998 * 14'd1631)) ^ (a ? 14'd11428 : 7256)) : 11403));
            
            4'd5: result_0337 = (14'd15895 << 2);
            
            4'd6: result_0337 = ((((~a) ^ ((14'd9597 ^ 14'd12380) ? (14'd13197 >> 1) : 4150)) + 14'd572) & ((14'd14245 >> 3) & 14'd11099));
            
            4'd7: result_0337 = (((((14'd339 << 3) | (a ? 14'd12770 : 14304)) - ((b * a) | (a ? 14'd971 : 10557))) << 2) * 14'd8492);
            
            4'd8: result_0337 = (((14'd5151 & a) - (b | (a | (b ^ b)))) ? 14'd1139 : 3779);
            
            4'd9: result_0337 = ((b | (~((14'd7449 + b) * (b + b)))) ^ (14'd12871 - (((a * 14'd7161) ^ (14'd1548 - b)) >> 3)));
            
            4'd10: result_0337 = ((((~b) | a) & (((14'd7061 >> 3) | (14'd16170 ? a : 16368)) + ((14'd14067 * 14'd9957) + (b * 14'd10190)))) - 14'd16375);
            
            4'd11: result_0337 = (14'd9266 * a);
            
            4'd12: result_0337 = (((((~14'd355) >> 1) + (a + b)) * b) & (14'd6985 + 14'd2346));
            
            4'd13: result_0337 = ((~(((14'd10708 * 14'd2534) >> 1) * 14'd6324)) << 3);
            
            default: result_0337 = 14'd11013;
        endcase
    end

endmodule
        