
module simple_alu_0477(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0477
);

    always @(*) begin
        case(op)
            
            4'd0: result_0477 = (((((14'd14125 - 14'd8180) >> 2) | ((b ^ 14'd16221) + (14'd11897 & 14'd10456))) + ((14'd13425 ^ 14'd494) ? (a * 14'd6628) : 11233)) + 14'd2629);
            
            4'd1: result_0477 = (b * (((14'd6691 * (14'd551 | 14'd12395)) * (14'd11571 ^ (14'd13855 - 14'd11254))) - (~14'd14206)));
            
            4'd2: result_0477 = (((~(14'd1021 + (14'd9243 >> 2))) << 3) ? a : 15901);
            
            4'd3: result_0477 = ((((14'd916 ^ 14'd570) << 1) - b) & 14'd10711);
            
            4'd4: result_0477 = (14'd5415 & (a << 2));
            
            4'd5: result_0477 = (((((14'd4377 + 14'd9662) ^ (14'd15331 * 14'd13878)) * 14'd6129) ^ ((14'd10168 ? (14'd15700 >> 3) : 3030) | ((14'd7209 ^ 14'd9460) + 14'd5113))) >> 2);
            
            4'd6: result_0477 = ((~(((14'd12223 | a) & b) << 2)) ? ((((~b) ? (b - a) : 3493) * a) << 3) : 15098);
            
            4'd7: result_0477 = (a << 2);
            
            4'd8: result_0477 = ((((14'd13360 ^ 14'd11218) << 1) << 1) >> 1);
            
            4'd9: result_0477 = (~14'd5468);
            
            4'd10: result_0477 = (((((a ? 14'd16059 : 1674) >> 3) ? b : 7933) ^ (b | ((b - 14'd5028) >> 1))) * (~14'd15811));
            
            4'd11: result_0477 = (14'd11986 * (b - (a + 14'd11339)));
            
            default: result_0477 = 14'd15055;
        endcase
    end

endmodule
        