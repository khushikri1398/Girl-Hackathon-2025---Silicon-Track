
module simple_alu_0272(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0272
);

    always @(*) begin
        case(op)
            
            4'd0: result_0272 = ((((14'd14559 ? (14'd3510 ^ b) : 11742) & ((a + 14'd12274) * (14'd9701 - 14'd11730))) & 14'd11686) ^ b);
            
            4'd1: result_0272 = (((((b ? 14'd1636 : 10105) - (a << 2)) - a) - (((14'd4033 >> 1) | (a ? a : 10029)) + ((14'd7488 * 14'd15833) >> 1))) | (~14'd11857));
            
            4'd2: result_0272 = ((a << 1) << 2);
            
            4'd3: result_0272 = (((~b) ^ (((b ^ 14'd8125) ^ (14'd1963 * b)) | (14'd8207 - 14'd1807))) - ((((14'd5300 * 14'd10177) + (14'd6236 - 14'd2295)) - ((14'd14039 - 14'd12199) * (14'd8841 << 2))) >> 2));
            
            4'd4: result_0272 = (14'd2394 >> 3);
            
            default: result_0272 = 14'd1009;
        endcase
    end

endmodule
        