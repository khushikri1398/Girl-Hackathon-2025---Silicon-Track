
module simple_alu_0162(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0162
);

    always @(*) begin
        case(op)
            
            4'd0: result_0162 = (a & (14'd11139 * 14'd14268));
            
            4'd1: result_0162 = (14'd15154 | ((~(14'd4739 + (14'd14339 ^ 14'd2458))) ? ((14'd13414 & (14'd8654 | a)) ? ((14'd12411 ^ 14'd14100) ^ (~14'd13276)) : 2234) : 10186));
            
            4'd2: result_0162 = (((~(a - 14'd5872)) >> 3) ? ((14'd9195 * ((14'd4431 ? b : 15183) ? (14'd4376 * 14'd5393) : 5651)) | (((b >> 1) << 3) ? 14'd7844 : 8514)) : 77);
            
            4'd3: result_0162 = (14'd2948 ^ ((((14'd5316 ? 14'd14414 : 8512) - (~a)) & b) ^ ((14'd6478 ^ 14'd6095) ? (b & 14'd5724) : 946)));
            
            4'd4: result_0162 = (((~a) - 14'd5533) * 14'd7559);
            
            4'd5: result_0162 = (~((a & ((14'd4307 >> 1) & (a * 14'd14236))) - b));
            
            4'd6: result_0162 = (14'd15858 >> 1);
            
            4'd7: result_0162 = (b ? (b & 14'd2779) : 10064);
            
            4'd8: result_0162 = (~(b >> 2));
            
            4'd9: result_0162 = ((b ? 14'd11111 : 7249) << 3);
            
            4'd10: result_0162 = (~(((~(14'd15371 << 1)) + ((a ^ 14'd2642) << 3)) ^ (14'd4640 * b)));
            
            4'd11: result_0162 = (((((14'd10002 >> 1) << 1) ^ (14'd9811 * (~a))) - (~((14'd9269 * a) & (14'd708 & 14'd10394)))) << 3);
            
            default: result_0162 = b;
        endcase
    end

endmodule
        