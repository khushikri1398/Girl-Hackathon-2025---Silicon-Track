
module simple_alu_0588(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0588
);

    always @(*) begin
        case(op)
            
            4'd0: result_0588 = (((14'd15711 + (14'd9901 ? 14'd15019 : 3855)) | ((14'd4384 ^ 14'd14557) >> 1)) ? ((((b & 14'd12234) << 2) * ((14'd6212 ^ 14'd7392) ? (14'd2402 >> 3) : 867)) << 3) : 10975);
            
            4'd1: result_0588 = (((((14'd3706 << 3) + (14'd8046 * a)) - a) >> 3) >> 1);
            
            4'd2: result_0588 = ((~14'd2396) * ((((14'd12124 * 14'd1218) << 1) + (14'd8072 | 14'd1746)) * ((14'd9623 | a) + ((14'd15744 ^ 14'd11768) ^ (14'd5882 | 14'd6252)))));
            
            4'd3: result_0588 = (b & (((14'd16005 ^ (a - 14'd14599)) * ((~14'd6922) & (~b))) * ((14'd8028 >> 3) + (~(14'd8834 ? a : 11231)))));
            
            4'd4: result_0588 = ((((14'd2571 << 1) << 1) | (((a * 14'd15013) ? b : 14838) - b)) >> 2);
            
            4'd5: result_0588 = (((((14'd13586 ? 14'd2686 : 8012) * 14'd14395) ? ((a ^ 14'd2679) | (14'd6428 + 14'd2271)) : 13720) << 3) ? ((b & ((a & 14'd6412) << 1)) ? (((b & 14'd538) ^ 14'd6364) & ((a - 14'd13913) - 14'd10131)) : 13436) : 4352);
            
            4'd6: result_0588 = (~14'd8686);
            
            4'd7: result_0588 = ((((~(14'd14649 - a)) >> 3) ^ (~14'd9388)) | ((b ^ 14'd6358) << 2));
            
            4'd8: result_0588 = ((((b & (14'd5010 - b)) - a) | b) << 2);
            
            4'd9: result_0588 = (((((14'd2803 << 2) & (b << 2)) + (~(a >> 3))) << 2) * ((a + a) & ((b << 3) ^ 14'd54)));
            
            4'd10: result_0588 = (((((14'd5540 << 1) >> 2) & 14'd11338) << 2) + ((((14'd12631 << 2) + (b ? 14'd742 : 14251)) >> 2) | (((14'd2795 + a) ? (a ? b : 15158) : 20) - (14'd116 * (14'd6484 | b)))));
            
            4'd11: result_0588 = (14'd2723 * 14'd16239);
            
            4'd12: result_0588 = (((~((a << 1) ? (14'd14983 & b) : 14621)) + (((a + 14'd4371) - a) * (~(14'd3416 ^ 14'd7544)))) & ((14'd6691 << 2) << 1));
            
            4'd13: result_0588 = (((b ^ ((a * 14'd627) >> 2)) ^ (((b ? 14'd5221 : 11687) ? (14'd12337 & a) : 9506) | ((14'd10824 << 3) ? (14'd12234 ^ 14'd12214) : 13151))) ^ (14'd2268 ^ a));
            
            default: result_0588 = 14'd460;
        endcase
    end

endmodule
        