
module simple_alu_0701(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0701
);

    always @(*) begin
        case(op)
            
            4'd0: result_0701 = (~((((b & 14'd15796) * (~a)) << 2) + 14'd8536));
            
            4'd1: result_0701 = (14'd9640 - (((a ^ (14'd8359 ^ 14'd14449)) + ((~14'd12265) * (14'd4602 - 14'd7403))) | b));
            
            4'd2: result_0701 = (((((14'd3783 * a) + (14'd4819 + 14'd10379)) >> 1) ? 14'd8903 : 9785) * (14'd9471 ? (~(~(b - 14'd5531))) : 6297));
            
            4'd3: result_0701 = (14'd10141 * (~((~(a >> 3)) ? (a - (~14'd5307)) : 3688)));
            
            4'd4: result_0701 = ((14'd2726 << 2) + (14'd3309 * (14'd15612 ? ((14'd11826 >> 1) & (14'd9823 * 14'd347)) : 13171)));
            
            4'd5: result_0701 = ((a >> 3) ? (~(((~14'd9232) - (14'd6457 >> 3)) * (14'd7318 ^ (14'd6388 + 14'd5025)))) : 1401);
            
            4'd6: result_0701 = (((((14'd6112 * 14'd2260) >> 1) - ((14'd10021 | a) & (b ^ 14'd1396))) ? a : 3342) - (~(14'd15919 & ((14'd15909 << 3) ? (14'd13690 >> 1) : 15697))));
            
            4'd7: result_0701 = ((14'd6431 ^ (14'd7136 | a)) ? ((((14'd14424 - b) + (14'd3520 & a)) << 2) >> 2) : 3992);
            
            4'd8: result_0701 = (14'd2987 ^ ((a * (14'd5122 | (14'd10477 ? 14'd12855 : 10571))) - ((14'd11542 ^ (14'd1611 ? 14'd4350 : 13648)) * a)));
            
            4'd9: result_0701 = ((b | (~((a << 3) ? 14'd2353 : 12823))) - ((((14'd7158 ? b : 8837) << 1) - ((14'd5482 & 14'd10556) * (14'd4429 >> 3))) << 3));
            
            default: result_0701 = 14'd2560;
        endcase
    end

endmodule
        