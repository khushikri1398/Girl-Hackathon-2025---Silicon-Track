
module simple_alu_0708(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0708
);

    always @(*) begin
        case(op)
            
            4'd0: result_0708 = ((~((b & (14'd5276 << 3)) << 2)) << 1);
            
            4'd1: result_0708 = (((b - b) & ((14'd4057 * a) >> 1)) + b);
            
            4'd2: result_0708 = (((((14'd6463 + b) + (14'd10662 ? a : 3150)) ^ ((a - 14'd14979) * (14'd14654 << 3))) - (((a & 14'd3049) ^ 14'd8215) | ((14'd6155 - 14'd1635) >> 1))) ? ((((a << 2) ? (14'd15388 + b) : 5617) ^ ((14'd14072 ? 14'd3340 : 13) ? 14'd8108 : 2138)) * (~(b | 14'd10933))) : 14509);
            
            4'd3: result_0708 = (((14'd1121 - ((14'd3081 >> 2) ? (14'd10713 & 14'd7079) : 14765)) ? ((14'd7859 ? (b - 14'd12270) : 427) & ((b >> 2) >> 3)) : 3362) & ((((14'd10863 & 14'd4664) ^ (14'd8133 >> 2)) << 2) | (14'd4405 ^ 14'd10630)));
            
            4'd4: result_0708 = (((((a + a) << 3) ? 14'd10647 : 8537) * (((b & 14'd9340) << 1) << 2)) - 14'd6439);
            
            4'd5: result_0708 = (~((14'd2257 & a) >> 3));
            
            4'd6: result_0708 = (14'd14606 ? (~(14'd5692 << 3)) : 14447);
            
            4'd7: result_0708 = (~14'd7916);
            
            4'd8: result_0708 = (((((b >> 3) ^ (~b)) * a) << 3) + (((14'd7774 + (14'd10607 >> 2)) | b) ? ((a * 14'd13001) * ((a + 14'd9431) + b)) : 8707));
            
            4'd9: result_0708 = (((((14'd916 * 14'd4841) | 14'd6721) * ((14'd13880 << 1) * (14'd5424 - 14'd11026))) ^ (((14'd10213 + b) >> 2) >> 3)) ^ ((14'd2830 | (14'd12635 ^ 14'd12168)) >> 2));
            
            4'd10: result_0708 = (((a << 2) | 14'd13264) << 2);
            
            4'd11: result_0708 = ((((14'd13519 & (a & b)) & a) | a) >> 3);
            
            4'd12: result_0708 = (((((~14'd10537) & (~b)) - (14'd14725 - b)) << 3) - ((((14'd4948 + b) ? (14'd13480 << 1) : 10276) | ((14'd15435 | a) + a)) & (((~14'd14381) ^ 14'd1046) >> 2)));
            
            4'd13: result_0708 = ((((~(14'd3195 ? 14'd10637 : 13402)) - 14'd14680) ^ b) << 1);
            
            4'd14: result_0708 = ((~(b - ((14'd14458 * 14'd16252) & (b >> 1)))) >> 2);
            
            4'd15: result_0708 = (((~((14'd12926 & 14'd13834) & (14'd12149 << 3))) + (((~14'd10970) & b) * ((b & 14'd11746) ? (a ^ 14'd12051) : 3709))) | ((14'd10589 + ((a | b) ^ (14'd9752 - 14'd15422))) - (((b | b) + 14'd1816) << 1)));
            
            default: result_0708 = 14'd6285;
        endcase
    end

endmodule
        