
module simple_alu_0807(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0807
);

    always @(*) begin
        case(op)
            
            4'd0: result_0807 = ((14'd12099 & (14'd3951 * ((14'd12076 & 14'd5892) << 1))) ? (~(((14'd15961 * a) & 14'd9598) & ((~a) << 1))) : 3430);
            
            4'd1: result_0807 = (((((~a) | (~14'd10725)) << 1) ^ (((14'd11061 | 14'd13039) | (a ^ 14'd15987)) << 1)) * ((((a | 14'd13265) * (b & 14'd11048)) ^ (14'd9907 >> 2)) + (((14'd5499 | 14'd15636) ^ (a >> 1)) ^ ((a - 14'd13275) ^ (14'd12654 ? 14'd14085 : 8560)))));
            
            4'd2: result_0807 = (((14'd10191 << 3) ^ 14'd12721) - (((14'd10445 & a) * ((b ^ 14'd12942) + b)) ^ (((14'd12279 >> 1) & (a ? a : 8261)) - 14'd5174)));
            
            4'd3: result_0807 = (((14'd10698 + (~a)) | (14'd16335 * ((14'd8052 - b) << 1))) ^ (14'd2066 + (((14'd9926 ^ 14'd9922) * (a | 14'd14718)) + ((14'd10592 ^ 14'd8819) + (b | b)))));
            
            4'd4: result_0807 = ((~14'd1901) * ((14'd12173 - b) & ((14'd11239 | 14'd248) + ((14'd7212 & 14'd16083) ? (a * 14'd14257) : 2498))));
            
            4'd5: result_0807 = (((((14'd15341 >> 1) | (14'd5269 ? a : 586)) + ((14'd10594 + 14'd462) >> 3)) & (((14'd10111 >> 1) | (a | 14'd3375)) & (a ^ (14'd4909 ? 14'd8576 : 5694)))) << 2);
            
            4'd6: result_0807 = ((14'd1349 >> 1) ^ 14'd8154);
            
            4'd7: result_0807 = (a * 14'd8991);
            
            4'd8: result_0807 = ((a * (((14'd1876 & 14'd1557) + (a ^ a)) | b)) & (14'd1676 ^ (((b ^ b) - (14'd15409 >> 3)) >> 2)));
            
            4'd9: result_0807 = ((~a) * a);
            
            4'd10: result_0807 = ((b + (14'd5425 << 3)) - (((14'd5021 ? (~14'd1687) : 8484) - ((14'd15903 | 14'd311) ? (b & a) : 5912)) << 3));
            
            4'd11: result_0807 = ((((14'd6880 << 2) >> 3) | b) ? ((((a | a) >> 1) << 3) << 1) : 1198);
            
            4'd12: result_0807 = (((~14'd15301) ^ (((14'd8669 + 14'd6663) | (b ? b : 1402)) * ((a + a) ^ (b - b)))) - 14'd6210);
            
            4'd13: result_0807 = (((~((14'd4419 | b) | (14'd3188 ? b : 1814))) & (~((14'd15318 * b) << 2))) ^ (14'd4443 & (14'd12692 - ((b - b) >> 2))));
            
            default: result_0807 = a;
        endcase
    end

endmodule
        