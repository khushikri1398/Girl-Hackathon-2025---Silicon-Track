
module simple_alu_0779(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0779
);

    always @(*) begin
        case(op)
            
            4'd0: result_0779 = (((a - ((a ^ 14'd12113) - (~a))) - (~(a ? (14'd12461 | 14'd9523) : 6578))) * (~(((14'd4922 << 1) << 2) & (~(14'd11911 >> 2)))));
            
            4'd1: result_0779 = (14'd4862 | ((((14'd6096 << 2) - (14'd14991 | 14'd15171)) ? (~(~b)) : 2352) ^ 14'd14717));
            
            4'd2: result_0779 = ((14'd15076 & (14'd10486 >> 2)) ? 14'd15413 : 8169);
            
            4'd3: result_0779 = (14'd3596 - (b - (((14'd4930 ^ 14'd6209) ^ 14'd13849) - (~a))));
            
            4'd4: result_0779 = (~14'd9837);
            
            4'd5: result_0779 = (b << 2);
            
            4'd6: result_0779 = (b ? ((((a - 14'd995) + (b >> 1)) | ((~a) ? 14'd10859 : 11423)) << 1) : 1662);
            
            4'd7: result_0779 = (14'd54 | (14'd8820 & b));
            
            default: result_0779 = 14'd12769;
        endcase
    end

endmodule
        