
module simple_alu_0409(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0409
);

    always @(*) begin
        case(op)
            
            4'd0: result_0409 = ((14'd11774 * 14'd10247) ? a : 8659);
            
            4'd1: result_0409 = (14'd1843 - (14'd6762 << 2));
            
            4'd2: result_0409 = (((((14'd5591 & 14'd8217) - b) ^ ((14'd1545 ? a : 14609) + (14'd2859 ^ 14'd6184))) & (a - 14'd3233)) | 14'd5528);
            
            4'd3: result_0409 = (((((a & 14'd10258) ? (14'd9881 >> 3) : 8911) ^ a) - ((a ? a : 14165) + (14'd12466 ? (b ? 14'd7287 : 6178) : 761))) ^ (((~14'd5094) | a) - 14'd2140));
            
            4'd4: result_0409 = (((((14'd7604 >> 3) - a) & ((b & 14'd10920) << 3)) - (~(14'd2339 & 14'd1607))) ^ ((~(~(14'd213 | 14'd6317))) | (~14'd3969)));
            
            4'd5: result_0409 = ((((a + (~14'd15590)) ^ 14'd1165) << 1) - (14'd8183 >> 2));
            
            4'd6: result_0409 = (~(b << 2));
            
            4'd7: result_0409 = (14'd5153 | (14'd10506 | (a ^ ((a & 14'd7937) | 14'd5292))));
            
            4'd8: result_0409 = (~14'd2458);
            
            4'd9: result_0409 = (((b ? ((14'd5405 * 14'd13224) & (a | b)) : 13934) ^ (14'd8290 & ((b ? a : 12731) | 14'd15982))) | (14'd1503 & 14'd10271));
            
            4'd10: result_0409 = ((~(((14'd13609 * a) ? (14'd7242 | 14'd8916) : 4759) ^ 14'd5161)) - a);
            
            4'd11: result_0409 = (((~(a ^ (b ^ b))) | 14'd5309) & (((14'd10188 << 1) >> 3) + (~14'd6705)));
            
            4'd12: result_0409 = (14'd15713 >> 3);
            
            4'd13: result_0409 = ((a >> 2) | (((a << 2) - ((~14'd1962) << 2)) & ((a * (~14'd13609)) ? 14'd12600 : 11022)));
            
            default: result_0409 = b;
        endcase
    end

endmodule
        