
module simple_alu_0814(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0814
);

    always @(*) begin
        case(op)
            
            4'd0: result_0814 = (a & ((14'd10391 * ((14'd1647 | a) | (a ? 14'd15370 : 6217))) ^ (((~a) ^ (14'd12520 | 14'd2934)) ? ((14'd15011 & 14'd12491) * (14'd1095 + a)) : 11198)));
            
            4'd1: result_0814 = ((((14'd1401 * 14'd6837) | ((b & 14'd8402) + (14'd16210 - 14'd2649))) ? ((14'd6475 * (b ^ 14'd6688)) + (~14'd6679)) : 5078) | 14'd6103);
            
            4'd2: result_0814 = (((b & (b - (14'd11836 + a))) << 1) >> 2);
            
            4'd3: result_0814 = (((~((b ^ 14'd6764) ^ (a >> 3))) | (b * (b ^ 14'd2161))) - (14'd3021 | (~14'd1910)));
            
            4'd4: result_0814 = (((((a - 14'd1712) + (a | 14'd6786)) & (a & (a ^ 14'd7184))) ^ 14'd7141) | ((((14'd15111 - a) ^ (14'd7963 | 14'd11989)) + 14'd12820) | ((14'd10283 << 2) & b)));
            
            4'd5: result_0814 = ((14'd11940 >> 2) ^ ((((b >> 3) + (14'd12736 << 1)) - a) >> 1));
            
            4'd6: result_0814 = (14'd2179 - 14'd10189);
            
            4'd7: result_0814 = (~b);
            
            4'd8: result_0814 = ((14'd9719 * b) ^ (((~(14'd3458 ^ 14'd9501)) - ((~14'd4134) >> 2)) & (~((a >> 2) & 14'd10992))));
            
            4'd9: result_0814 = ((14'd10081 + (14'd5502 - ((a + 14'd2137) >> 2))) | (14'd6873 & (14'd13298 ^ (~(14'd11882 - 14'd12151)))));
            
            4'd10: result_0814 = (14'd5783 ? 14'd7147 : 12145);
            
            4'd11: result_0814 = (((((b | 14'd10901) >> 1) ^ ((14'd731 ^ a) >> 1)) - ((~14'd2654) << 1)) << 3);
            
            4'd12: result_0814 = ((b >> 3) * (14'd583 & 14'd15631));
            
            default: result_0814 = b;
        endcase
    end

endmodule
        