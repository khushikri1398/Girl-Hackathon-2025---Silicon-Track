
module simple_alu_0377(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0377
);

    always @(*) begin
        case(op)
            
            4'd0: result_0377 = ((b & 14'd2647) ^ (14'd4218 + (((a + b) - (b >> 1)) + (b ? a : 8850))));
            
            4'd1: result_0377 = ((a << 3) & 14'd7254);
            
            4'd2: result_0377 = (14'd11940 * ((((14'd7768 * b) & (14'd11511 ? a : 2376)) ? ((b ? 14'd11632 : 15392) << 1) : 8565) & ((~14'd6265) + 14'd13435)));
            
            4'd3: result_0377 = (~(14'd801 - 14'd4276));
            
            4'd4: result_0377 = (((14'd12416 & (14'd8349 - 14'd16338)) | (~14'd10695)) * ((~((14'd991 & 14'd2551) | (14'd2068 << 2))) * (b - 14'd5746)));
            
            4'd5: result_0377 = ((14'd13067 << 3) * 14'd9767);
            
            4'd6: result_0377 = ((((14'd15081 * (b * 14'd9832)) - b) & (14'd7962 >> 3)) & 14'd10386);
            
            4'd7: result_0377 = (((~(~(14'd2544 >> 1))) - ((14'd15985 & (14'd8042 & 14'd4891)) << 1)) - 14'd1633);
            
            4'd8: result_0377 = (~((((14'd7952 * 14'd14344) ^ 14'd22) ? 14'd7318 : 16370) >> 2));
            
            4'd9: result_0377 = (((a - a) * (((14'd1177 << 1) >> 3) - ((a & b) ^ (~a)))) >> 3);
            
            default: result_0377 = a;
        endcase
    end

endmodule
        