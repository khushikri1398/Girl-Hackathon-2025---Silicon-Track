
module simple_alu_0998(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0998
);

    always @(*) begin
        case(op)
            
            4'd0: result_0998 = ((a ? (((~14'd13353) - (~14'd8079)) << 1) : 430) & a);
            
            4'd1: result_0998 = (((((b << 2) ? (~14'd1909) : 8411) >> 3) * (((a << 1) + (14'd1820 >> 3)) >> 1)) ? 14'd15939 : 16116);
            
            4'd2: result_0998 = (((b - ((a ^ a) ^ (14'd9662 & a))) | (((b * 14'd1656) + (b ^ 14'd15886)) ^ 14'd15053)) * (14'd160 - 14'd4994));
            
            4'd3: result_0998 = (14'd8045 + a);
            
            4'd4: result_0998 = ((14'd11135 * b) - ((((14'd2534 ? 14'd14930 : 119) - 14'd2982) >> 1) ^ (((14'd5063 ^ 14'd15742) >> 2) & 14'd11329)));
            
            4'd5: result_0998 = ((~(b * 14'd11261)) & ((14'd15663 - 14'd188) & (~(14'd14006 ^ (14'd2445 ? 14'd6803 : 13834)))));
            
            4'd6: result_0998 = ((14'd13635 ? a : 3766) + ((((b << 3) & 14'd757) >> 3) & ((a + (b << 1)) << 2)));
            
            4'd7: result_0998 = (14'd14255 & 14'd11714);
            
            4'd8: result_0998 = (14'd10665 ? (a << 1) : 4155);
            
            4'd9: result_0998 = ((((14'd8877 * (14'd12979 | 14'd14691)) ? ((~14'd7946) - (a | 14'd7213)) : 2889) + (((a ? b : 11517) + (~14'd10584)) << 1)) * (14'd2764 | (((b ? 14'd2528 : 5094) << 1) | ((14'd3744 >> 3) | (~14'd7546)))));
            
            4'd10: result_0998 = (((14'd15714 ? b : 13697) >> 1) >> 2);
            
            4'd11: result_0998 = (~((14'd2075 - b) * (((14'd3196 | 14'd4626) - (a & b)) * (~(14'd3921 ? 14'd14432 : 13590)))));
            
            4'd12: result_0998 = (14'd3403 - a);
            
            4'd13: result_0998 = (14'd4992 - (((14'd12348 - 14'd14038) + (~b)) * (((14'd4319 * 14'd464) & (b >> 1)) >> 3)));
            
            default: result_0998 = 14'd3286;
        endcase
    end

endmodule
        