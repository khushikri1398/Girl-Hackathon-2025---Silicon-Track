
module simple_alu_0536(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0536
);

    always @(*) begin
        case(op)
            
            4'd0: result_0536 = ((((~(14'd8443 << 1)) * 14'd3372) + (~(14'd7182 << 2))) << 1);
            
            4'd1: result_0536 = (~(a ^ (14'd2391 + ((a ^ a) - (14'd2141 ? 14'd5754 : 8130)))));
            
            4'd2: result_0536 = (((~(b * (14'd14621 - 14'd8934))) ? (~14'd865) : 9267) - ((a * (14'd3925 ^ (a ^ a))) ? (((14'd5009 - 14'd4976) | (14'd6607 ^ 14'd10612)) ? 14'd14466 : 13376) : 5117));
            
            4'd3: result_0536 = ((14'd15839 << 2) * (14'd11361 & (((14'd8594 ^ 14'd9013) << 2) >> 1)));
            
            4'd4: result_0536 = (((((b * a) + (14'd1179 - 14'd2536)) << 2) >> 2) ^ 14'd1607);
            
            4'd5: result_0536 = (((((14'd14255 ^ 14'd9057) ^ 14'd5012) ? a : 13705) ^ (14'd15421 + ((14'd3894 ^ 14'd12262) * (a | b)))) | ((14'd120 >> 1) | (14'd5277 >> 3)));
            
            4'd6: result_0536 = (14'd13758 * 14'd6803);
            
            4'd7: result_0536 = ((14'd4278 * (14'd2431 & ((14'd6118 << 3) & (14'd12971 + a)))) - (14'd8373 << 3));
            
            4'd8: result_0536 = ((((b ^ (14'd4332 & a)) ? (14'd11646 ^ (a | 14'd7253)) : 7808) ? (((14'd105 ^ 14'd7086) ? (14'd8179 & 14'd1045) : 12134) | 14'd907) : 1156) ^ (14'd7883 - (((14'd5579 - 14'd8224) << 3) >> 3)));
            
            4'd9: result_0536 = (((((a ? 14'd6296 : 13954) >> 2) - ((~b) ? (14'd5085 & 14'd1029) : 5308)) >> 2) >> 2);
            
            4'd10: result_0536 = ((14'd15514 * (((~14'd15816) ? (b | b) : 7986) ^ ((14'd15280 | 14'd7931) + (14'd2351 - 14'd9621)))) | a);
            
            4'd11: result_0536 = (14'd2040 * ((((14'd1663 & 14'd9836) ^ (14'd15844 + 14'd15102)) | b) << 1));
            
            4'd12: result_0536 = (b ^ ((((a << 2) * (~b)) ? ((14'd3940 & a) * b) : 15282) - (((b & b) ? (~14'd14944) : 10522) << 1)));
            
            4'd13: result_0536 = (~((((b & a) | (b ^ 14'd13970)) ^ 14'd15531) >> 1));
            
            default: result_0536 = b;
        endcase
    end

endmodule
        