
module simple_alu_0288(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0288
);

    always @(*) begin
        case(op)
            
            4'd0: result_0288 = ((a << 2) >> 3);
            
            4'd1: result_0288 = (a >> 3);
            
            4'd2: result_0288 = (a + ((((14'd9605 | a) ^ (b + 14'd159)) ? ((a + a) & (14'd10597 & b)) : 2593) - ((~(14'd11493 << 1)) * ((14'd4657 & 14'd14986) ? (b >> 1) : 16311))));
            
            4'd3: result_0288 = (((((14'd16273 ? 14'd3622 : 2123) & (a * 14'd3097)) * b) | (((~14'd12937) | (14'd3132 ? 14'd5506 : 10763)) << 2)) | ((b * 14'd2243) & 14'd12210));
            
            4'd4: result_0288 = ((((14'd14559 + (14'd3780 - b)) ? 14'd4781 : 11995) & ((b & (14'd1975 + 14'd1404)) - (~(14'd6402 ? b : 477)))) & (b | ((~(14'd15535 >> 2)) * ((~14'd8122) << 1))));
            
            4'd5: result_0288 = ((b * (a + (14'd5542 << 1))) - a);
            
            4'd6: result_0288 = ((14'd5717 | (14'd10138 >> 1)) - (14'd943 ^ (((b * b) ? (b | b) : 3462) & ((b - b) | 14'd14998))));
            
            4'd7: result_0288 = (((((14'd6572 ^ 14'd15193) * (14'd11174 ? a : 894)) * 14'd5030) ^ (a & ((14'd15496 | 14'd6117) ^ a))) ? ((14'd9623 & ((b | 14'd11764) | (a ? b : 13406))) + (((14'd1791 - 14'd2260) - (14'd10073 ? 14'd8058 : 12513)) | ((14'd5886 ^ 14'd4818) | (14'd5045 | b)))) : 15507);
            
            4'd8: result_0288 = (((b & ((~b) ^ (14'd7289 | a))) & ((~b) - ((a | 14'd1412) << 3))) - (~(~((a ? 14'd4118 : 4086) ? (14'd16352 * a) : 13376))));
            
            4'd9: result_0288 = (14'd8342 - b);
            
            4'd10: result_0288 = ((b & (((14'd435 & a) | a) & 14'd12076)) + (14'd10261 + a));
            
            default: result_0288 = b;
        endcase
    end

endmodule
        