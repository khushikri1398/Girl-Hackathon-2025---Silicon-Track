
module simple_alu_0360(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0360
);

    always @(*) begin
        case(op)
            
            4'd0: result_0360 = (14'd3006 & (14'd12587 ? (((b ^ 14'd6335) + 14'd13963) ? 14'd4553 : 746) : 13694));
            
            4'd1: result_0360 = ((((14'd3324 + (a ? a : 12007)) * ((14'd8481 ^ 14'd12558) ? (a + 14'd15500) : 10850)) | (((b & a) >> 1) - ((a - b) - (~a)))) | a);
            
            4'd2: result_0360 = ((((a & (14'd12001 ? 14'd14186 : 6684)) & (14'd1461 + (b & 14'd13888))) | (((~a) | (b + 14'd10175)) * ((14'd14360 & 14'd4084) & (b & b)))) ? b : 13883);
            
            4'd3: result_0360 = ((((14'd13811 - (a - 14'd3514)) | 14'd2657) | (b ^ ((14'd9855 & a) >> 2))) | ((((~14'd16170) << 2) & 14'd7175) ? ((~(14'd8755 + 14'd16282)) ^ ((b + a) >> 1)) : 14320));
            
            4'd4: result_0360 = (b + a);
            
            4'd5: result_0360 = ((((~a) ? ((14'd2160 ^ b) ? (14'd3816 & 14'd7064) : 6240) : 3543) >> 2) * 14'd4999);
            
            4'd6: result_0360 = (((~((~a) - (14'd6834 + 14'd6185))) - (((14'd9897 & b) & 14'd2353) >> 2)) + ((((b << 3) - 14'd9788) << 3) + b));
            
            default: result_0360 = b;
        endcase
    end

endmodule
        