
module simple_alu_0451(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0451
);

    always @(*) begin
        case(op)
            
            4'd0: result_0451 = (((14'd3366 >> 2) & (14'd2444 ? ((14'd14914 * 14'd14106) >> 1) : 6052)) >> 2);
            
            4'd1: result_0451 = (a ? 14'd15113 : 10066);
            
            4'd2: result_0451 = ((14'd519 - (~a)) << 2);
            
            4'd3: result_0451 = (((((14'd3008 ? 14'd3647 : 8724) >> 2) ^ ((14'd329 + 14'd11660) | (b - 14'd8126))) & (a ^ ((14'd10506 | b) >> 3))) >> 1);
            
            4'd4: result_0451 = (((~(~(14'd9337 | a))) & (b - ((a & b) - (14'd926 & 14'd4118)))) << 3);
            
            4'd5: result_0451 = (((((14'd2159 & 14'd8739) - (~14'd10420)) << 2) ^ (((14'd16198 | 14'd15129) | 14'd7146) ? (14'd5392 ? (14'd15081 - b) : 8611) : 4760)) | 14'd8242);
            
            4'd6: result_0451 = (((b | 14'd12343) | ((14'd10160 + (b - a)) + (b - (14'd5222 ? b : 15851)))) >> 1);
            
            4'd7: result_0451 = (((((b ^ b) | (14'd515 | 14'd3217)) & (14'd10908 & (a * 14'd9711))) >> 1) & ((~((14'd11115 | b) ? (~a) : 2403)) << 1));
            
            4'd8: result_0451 = (((~14'd8759) << 1) ? ((((b << 2) * (b * 14'd16187)) << 1) - ((14'd4976 + (b ^ 14'd5869)) ^ ((14'd13263 & 14'd2268) ^ (b << 2)))) : 108);
            
            4'd9: result_0451 = (((((~b) - (14'd12029 + b)) + ((14'd12633 + 14'd3404) - (b >> 1))) + 14'd15249) << 2);
            
            4'd10: result_0451 = (((14'd16039 - ((b ^ 14'd1512) * (a & 14'd16304))) | (((14'd8917 ^ b) - (14'd6629 & b)) ^ ((14'd10476 & a) ^ (a + a)))) - (((~(b ^ 14'd6659)) << 3) & (14'd187 ^ (14'd6898 ^ (a | 14'd9152)))));
            
            4'd11: result_0451 = ((((~14'd8574) - (14'd7646 | (~14'd5992))) << 3) | (14'd9212 * ((~a) << 3)));
            
            4'd12: result_0451 = (~((((~14'd2355) >> 1) - ((14'd16074 | b) * (14'd12137 & a))) ? (14'd15977 & ((14'd10117 ? 14'd14378 : 8982) ^ 14'd8769)) : 12822));
            
            4'd13: result_0451 = ((((a << 1) >> 3) ^ (((a ^ 14'd12735) | (a ^ b)) - ((a >> 2) * b))) << 3);
            
            default: result_0451 = 14'd9573;
        endcase
    end

endmodule
        