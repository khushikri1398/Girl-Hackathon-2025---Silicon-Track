
module simple_alu_0812(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0812
);

    always @(*) begin
        case(op)
            
            4'd0: result_0812 = (~(((~(~b)) >> 2) * ((~(14'd1144 >> 3)) + 14'd587)));
            
            4'd1: result_0812 = (((14'd7249 << 1) >> 1) * (a + (14'd2986 - b)));
            
            4'd2: result_0812 = (b & ((((a ? 14'd1195 : 4031) >> 3) << 3) - (b - 14'd15748)));
            
            4'd3: result_0812 = ((~(((b & 14'd5162) & 14'd14418) + b)) & a);
            
            4'd4: result_0812 = (~14'd12105);
            
            4'd5: result_0812 = (14'd2173 & (14'd8874 - 14'd3112));
            
            4'd6: result_0812 = (~((a - 14'd15219) << 3));
            
            4'd7: result_0812 = (((((b * 14'd10225) & (14'd15189 ^ 14'd10022)) & (~(14'd12707 | 14'd13595))) ? (((a | 14'd112) ? 14'd2547 : 2585) | ((b + b) | (~14'd16209))) : 12985) | (14'd2078 | 14'd6200));
            
            4'd8: result_0812 = (14'd11371 | (b * (14'd2988 | b)));
            
            4'd9: result_0812 = (b >> 1);
            
            4'd10: result_0812 = ((~(((14'd13905 >> 3) | (14'd10112 * 14'd12496)) ? (b ? (b & 14'd12707) : 2785) : 10191)) ^ 14'd6146);
            
            4'd11: result_0812 = ((b ? (((b ? 14'd14715 : 12274) | (b - a)) + ((~14'd8168) + (~b))) : 7255) + b);
            
            4'd12: result_0812 = (~14'd8318);
            
            4'd13: result_0812 = ((((14'd16219 ^ (~14'd14682)) >> 1) ^ ((14'd14023 * (14'd14020 << 2)) + a)) * ((14'd5888 - ((14'd5279 >> 3) ^ a)) + ((14'd10159 ? (b ? a : 495) : 8270) + ((14'd38 << 3) >> 2))));
            
            4'd14: result_0812 = (((((14'd9878 ? 14'd15610 : 14530) >> 1) ^ 14'd5348) >> 1) >> 1);
            
            default: result_0812 = a;
        endcase
    end

endmodule
        