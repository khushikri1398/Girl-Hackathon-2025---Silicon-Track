
module simple_alu_0383(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0383
);

    always @(*) begin
        case(op)
            
            4'd0: result_0383 = (b ? ((((14'd9170 + a) * (b ? b : 876)) - (14'd12922 >> 3)) * (((a + b) >> 1) * (14'd5574 + (14'd2180 + 14'd369)))) : 212);
            
            4'd1: result_0383 = (((((~14'd13892) * (a * 14'd4025)) - ((14'd14235 * b) & (14'd14520 - b))) ? 14'd11039 : 2494) >> 3);
            
            4'd2: result_0383 = (~(14'd16301 >> 2));
            
            4'd3: result_0383 = (((a * 14'd5816) ^ (b << 3)) - (((~(a * 14'd449)) ? (a ^ 14'd4415) : 9295) * 14'd3328));
            
            4'd4: result_0383 = (((((14'd1819 ^ 14'd639) >> 2) | 14'd7683) << 3) << 1);
            
            4'd5: result_0383 = ((b & (((b & a) - (14'd8657 ^ a)) << 1)) ^ ((a >> 3) ^ (~((~14'd13747) >> 3))));
            
            4'd6: result_0383 = (((((a + 14'd11309) << 1) ? ((~b) * (~14'd13515)) : 11467) << 1) * (((b & b) * (b * (14'd8399 ^ b))) ? (((a >> 1) << 1) ^ (14'd8431 + 14'd7739)) : 7429));
            
            4'd7: result_0383 = (((14'd6956 >> 1) + 14'd9856) * (((14'd3578 ? (~14'd1855) : 594) * ((14'd4923 << 3) | 14'd12545)) & 14'd15276));
            
            4'd8: result_0383 = (14'd11849 + ((14'd9524 | 14'd2430) ? (((14'd4720 << 3) >> 2) & 14'd6107) : 466));
            
            4'd9: result_0383 = (b - a);
            
            4'd10: result_0383 = (((~((14'd2713 * b) + (14'd15947 + 14'd15571))) | 14'd858) - 14'd4391);
            
            4'd11: result_0383 = (14'd8309 - (a & (14'd335 & (~(a ^ 14'd11018)))));
            
            4'd12: result_0383 = (((14'd9409 | (14'd13681 * b)) - a) + a);
            
            4'd13: result_0383 = (14'd6062 * ((((a + 14'd7024) + (a ^ 14'd4804)) >> 3) | (a ^ ((~a) | 14'd7038))));
            
            default: result_0383 = 14'd4719;
        endcase
    end

endmodule
        