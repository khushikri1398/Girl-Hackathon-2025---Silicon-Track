
module simple_alu_0221(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0221
);

    always @(*) begin
        case(op)
            
            4'd0: result_0221 = (((14'd4260 * (~(14'd8606 + a))) << 3) | (a * (((14'd4665 ^ a) | (14'd12955 ^ 14'd9353)) - ((~14'd5254) - (b + a)))));
            
            4'd1: result_0221 = (((((14'd10538 * 14'd13320) ^ 14'd4975) - ((14'd6092 * 14'd7453) - (14'd9606 + 14'd13923))) - 14'd3379) >> 1);
            
            4'd2: result_0221 = ((((14'd3071 * (14'd14752 * 14'd2470)) & ((14'd3624 >> 2) * (a << 2))) - 14'd55) ? (~14'd8684) : 9831);
            
            4'd3: result_0221 = ((((14'd10572 | (a * a)) * ((a & b) << 1)) | ((~14'd11438) << 2)) ? (14'd6319 << 3) : 16260);
            
            4'd4: result_0221 = (14'd948 + ((((14'd3255 - 14'd10091) << 3) >> 2) ^ ((14'd329 ^ (~14'd8135)) ^ b)));
            
            4'd5: result_0221 = (~(14'd2484 + ((a << 3) << 1)));
            
            4'd6: result_0221 = ((14'd6731 << 1) << 1);
            
            4'd7: result_0221 = ((b + (((a ? a : 8308) | (14'd14569 & 14'd15855)) * ((14'd3623 ^ 14'd3117) | 14'd8005))) >> 2);
            
            4'd8: result_0221 = ((14'd12878 | (((14'd1385 + b) - (a & 14'd13723)) >> 3)) * ((((b >> 1) ? (14'd13996 * 14'd6791) : 6397) << 3) | (((14'd3114 << 3) << 2) & ((b - a) << 3))));
            
            4'd9: result_0221 = ((((b - 14'd4772) >> 3) ^ (((b + 14'd3917) >> 2) >> 2)) - 14'd4957);
            
            4'd10: result_0221 = ((~14'd15412) << 1);
            
            4'd11: result_0221 = ((14'd14737 & b) - (((~14'd12422) + ((a ^ 14'd9623) >> 2)) & (((~b) * (a - 14'd4820)) + a)));
            
            4'd12: result_0221 = (~((((14'd5823 & 14'd2312) - 14'd6970) * b) | (((a | 14'd6433) + (14'd12166 >> 1)) >> 3)));
            
            default: result_0221 = a;
        endcase
    end

endmodule
        