
module simple_alu_0818(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0818
);

    always @(*) begin
        case(op)
            
            4'd0: result_0818 = (a >> 3);
            
            4'd1: result_0818 = (14'd13139 << 2);
            
            4'd2: result_0818 = (((~b) * b) + (b * (((14'd6815 | a) << 3) ? (14'd5185 ? (14'd10124 & 14'd4175) : 3659) : 10526)));
            
            4'd3: result_0818 = (((14'd9080 | ((14'd6944 ^ 14'd16237) >> 3)) * (((14'd6731 - b) | (b - a)) ^ 14'd9213)) - ((~((14'd5021 & b) << 2)) + (14'd7832 * 14'd13742)));
            
            4'd4: result_0818 = (~14'd15573);
            
            4'd5: result_0818 = (((14'd12286 << 1) | 14'd8227) | 14'd13596);
            
            4'd6: result_0818 = (a ? ((((14'd13700 | a) * (a + a)) << 1) ? (((14'd3411 + b) - (14'd2628 >> 3)) << 3) : 3007) : 8481);
            
            4'd7: result_0818 = (((((14'd3962 | a) * (b + 14'd1923)) | ((14'd4641 - 14'd666) ? 14'd1030 : 1516)) | (b ^ 14'd5866)) * (((~(14'd9548 ^ b)) & (~(b - a))) | (~(b & a))));
            
            4'd8: result_0818 = (((~((14'd12231 << 1) - (b ? a : 12026))) ? 14'd12119 : 637) ^ (b | (((14'd15174 * a) >> 1) ? ((a >> 1) * (14'd11552 << 1)) : 827)));
            
            4'd9: result_0818 = (~b);
            
            4'd10: result_0818 = ((14'd3615 | (14'd1970 * ((b >> 3) >> 1))) >> 1);
            
            4'd11: result_0818 = (b >> 3);
            
            4'd12: result_0818 = (a - (((~b) - 14'd4095) << 3));
            
            default: result_0818 = a;
        endcase
    end

endmodule
        