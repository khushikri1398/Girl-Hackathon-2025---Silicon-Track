
module simple_alu_0444(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0444
);

    always @(*) begin
        case(op)
            
            4'd0: result_0444 = (((((a - 14'd11696) + 14'd9708) << 1) ? (((b + 14'd7831) - 14'd8949) << 2) : 428) + (~(((b * 14'd11982) << 2) ? 14'd7465 : 2777)));
            
            4'd1: result_0444 = (a ? ((14'd15301 ? a : 2886) << 1) : 10094);
            
            4'd2: result_0444 = (((((b << 1) + (14'd3219 ? b : 16079)) >> 1) * (((14'd1339 << 1) ^ (~14'd6338)) ^ (14'd4772 ? (a * 14'd14463) : 12929))) ^ ((a ? ((a ^ a) + (14'd11918 >> 3)) : 14764) << 2));
            
            4'd3: result_0444 = (14'd10740 ? ((((14'd1348 ? 14'd11208 : 1540) | (14'd4396 + 14'd10486)) >> 2) + 14'd15715) : 587);
            
            4'd4: result_0444 = (((14'd5896 - a) * (((14'd14926 * a) | (a * 14'd2458)) ? 14'd14694 : 4603)) - (14'd13054 << 3));
            
            4'd5: result_0444 = (b << 3);
            
            4'd6: result_0444 = (14'd6699 ^ (a ? 14'd4626 : 8329));
            
            4'd7: result_0444 = (14'd16108 + 14'd8079);
            
            4'd8: result_0444 = (14'd4164 + (14'd4644 * 14'd7923));
            
            4'd9: result_0444 = ((((~(14'd9058 & 14'd5541)) | ((b ^ b) * (14'd12594 * 14'd8614))) ? (((~14'd12698) ^ (a * 14'd10500)) + ((a ? 14'd10226 : 10400) & (14'd15012 - b))) : 9457) ? (a ? ((14'd2239 - (14'd3607 ^ 14'd12333)) + 14'd15661) : 12411) : 11958);
            
            4'd10: result_0444 = (a >> 3);
            
            4'd11: result_0444 = (~((b - (14'd5205 >> 1)) & (((a * b) & 14'd9622) << 2)));
            
            4'd12: result_0444 = (14'd6513 * (14'd1753 | ((~(14'd4412 ? 14'd7935 : 4847)) >> 1)));
            
            default: result_0444 = 14'd14156;
        endcase
    end

endmodule
        