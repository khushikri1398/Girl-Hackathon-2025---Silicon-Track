
module simple_alu_0556(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0556
);

    always @(*) begin
        case(op)
            
            4'd0: result_0556 = (((((14'd38 + a) << 2) * 14'd16002) ? (14'd7357 + b) : 13470) + (b + 14'd369));
            
            4'd1: result_0556 = (14'd5673 & a);
            
            4'd2: result_0556 = ((((14'd5550 ^ (14'd12749 | 14'd2004)) & ((14'd15201 + 14'd7600) | (a | 14'd6027))) >> 2) | a);
            
            4'd3: result_0556 = ((a - 14'd4737) ^ ((((14'd6923 ? a : 14421) ? (14'd4861 | 14'd5445) : 875) << 2) & (~((14'd12014 & 14'd13793) ? (14'd15437 ^ 14'd4808) : 11640))));
            
            4'd4: result_0556 = (~((((a + 14'd1516) ^ 14'd14309) << 3) - (14'd2068 * ((~14'd6764) ? (14'd13442 ? 14'd9495 : 13227) : 13005))));
            
            4'd5: result_0556 = ((b ? (14'd508 * ((14'd12918 | a) * (14'd10929 >> 1))) : 11941) & ((((a - 14'd5876) & (14'd2063 ? b : 9395)) >> 1) ^ (((a << 3) ^ (~b)) ? ((a - 14'd1346) << 3) : 8215)));
            
            4'd6: result_0556 = ((((14'd11804 ^ (b >> 1)) - (14'd2723 & 14'd10017)) << 3) + ((14'd7201 | ((14'd8455 | 14'd6116) & (14'd8144 + b))) + ((~b) * ((14'd13836 - b) ? (14'd12420 ? 14'd11239 : 6261) : 15154))));
            
            4'd7: result_0556 = (14'd1859 * b);
            
            4'd8: result_0556 = ((14'd5121 ? ((a ^ (14'd6302 | b)) - 14'd15361) : 9421) ? (((a | (b << 1)) >> 1) - (14'd12214 - a)) : 12349);
            
            4'd9: result_0556 = (14'd15990 + ((((14'd14500 * b) | (a & a)) << 3) >> 1));
            
            4'd10: result_0556 = (((((b << 1) + 14'd1606) ^ (b ? (a << 1) : 3849)) & ((a * (b ? a : 13444)) + ((a - a) ^ b))) >> 1);
            
            4'd11: result_0556 = (14'd902 >> 1);
            
            4'd12: result_0556 = (14'd11581 >> 2);
            
            4'd13: result_0556 = (~((((14'd8053 + a) - (b + b)) * 14'd2510) - (~(~(b - 14'd14523)))));
            
            4'd14: result_0556 = ((b >> 3) + 14'd13159);
            
            default: result_0556 = b;
        endcase
    end

endmodule
        