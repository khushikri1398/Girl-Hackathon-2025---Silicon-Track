
module simple_alu_0009(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0009
);

    always @(*) begin
        case(op)
            
            4'd0: result_0009 = ((((14'd15689 | (14'd8041 * a)) & (14'd1993 ^ (a ? b : 3189))) + ((a * (a ^ 14'd9886)) * (b ? (b ^ b) : 7116))) * (14'd4622 >> 2));
            
            4'd1: result_0009 = (b ? ((((~14'd1599) & (14'd1204 * 14'd1423)) * ((~14'd3016) | (b + 14'd6059))) + (((a ? 14'd10739 : 2664) >> 2) & ((14'd13787 | 14'd8550) ? (14'd10203 & a) : 8206))) : 9377);
            
            4'd2: result_0009 = (14'd6114 * (((14'd11075 ^ 14'd7402) - ((a >> 1) ^ (14'd8109 >> 2))) - ((~(14'd15059 & b)) ^ ((b << 1) ? (~b) : 13109))));
            
            default: result_0009 = 14'd8378;
        endcase
    end

endmodule
        