
module simple_alu_0137(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0137
);

    always @(*) begin
        case(op)
            
            4'd0: result_0137 = (((((a - 14'd11713) & (14'd2810 * a)) >> 1) ? ((a >> 2) - ((14'd6301 & b) - 14'd12812)) : 11187) & (a - (((14'd11740 ? b : 16315) << 2) << 2)));
            
            4'd1: result_0137 = (a + (~((~(14'd9041 ^ 14'd5963)) << 1)));
            
            4'd2: result_0137 = ((a << 1) ? a : 9418);
            
            4'd3: result_0137 = ((((a & (14'd280 >> 3)) | 14'd87) & 14'd9062) | ((a * 14'd13423) ^ b));
            
            4'd4: result_0137 = (14'd4744 >> 2);
            
            4'd5: result_0137 = ((14'd15803 ? 14'd8653 : 9334) & ((14'd5235 * ((a * a) - 14'd11477)) | ((14'd16130 >> 3) & 14'd11976)));
            
            4'd6: result_0137 = ((~(((14'd16239 >> 2) - (a & 14'd14783)) + ((14'd1342 * 14'd14839) & (b | b)))) ? (~(a >> 2)) : 12434);
            
            4'd7: result_0137 = ((((14'd9031 + 14'd8026) + ((14'd8085 - b) | b)) << 2) ? (a << 3) : 5453);
            
            4'd8: result_0137 = (~(~(((b << 1) | a) * ((14'd24 ? 14'd2156 : 15916) << 1))));
            
            4'd9: result_0137 = (((((14'd2778 << 2) | 14'd776) ^ (a << 2)) ^ ((14'd13861 & (b >> 1)) * (a - (b >> 1)))) | ((~(14'd4665 * (14'd5292 - 14'd13556))) | (a - ((14'd8063 ? 14'd5441 : 2289) + (14'd7418 ? 14'd14162 : 15014)))));
            
            4'd10: result_0137 = (((14'd15107 ? (14'd15390 << 2) : 433) * (((14'd12666 | 14'd5673) << 2) ^ (a >> 2))) * ((((14'd14649 >> 1) << 2) | a) + (((b * 14'd13938) - (14'd10047 & 14'd13590)) * a)));
            
            4'd11: result_0137 = (14'd4742 ? 14'd261 : 15752);
            
            4'd12: result_0137 = (~((((a >> 3) | 14'd16133) ^ b) * a));
            
            default: result_0137 = b;
        endcase
    end

endmodule
        