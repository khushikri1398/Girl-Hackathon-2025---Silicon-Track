
module simple_alu_0949(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0949
);

    always @(*) begin
        case(op)
            
            4'd0: result_0949 = (((~14'd14632) ? (((a & a) ^ (b * 14'd5151)) * ((14'd7034 ^ b) >> 2)) : 8362) >> 1);
            
            4'd1: result_0949 = (~((14'd7789 - (14'd10497 + (14'd5541 | a))) >> 2));
            
            4'd2: result_0949 = ((~(((a ^ b) | a) - ((b | 14'd6875) ^ 14'd9518))) - ((14'd11047 * (~(14'd13669 ^ 14'd3147))) - (((14'd16144 << 3) * a) * 14'd13168)));
            
            4'd3: result_0949 = ((((~(14'd7870 ^ a)) | ((a - 14'd1947) >> 2)) & ((14'd5722 << 3) * ((14'd4860 * b) * (14'd8852 & b)))) | (~(14'd232 << 2)));
            
            4'd4: result_0949 = (14'd8666 ? (~14'd5279) : 14723);
            
            4'd5: result_0949 = (((((a & 14'd6350) + (a & 14'd13166)) ^ ((14'd1987 ? 14'd838 : 5186) | (14'd2915 ? b : 2386))) << 2) - ((((b ? a : 4469) + b) * (b & b)) & (a & 14'd13128)));
            
            4'd6: result_0949 = (14'd5225 + (14'd1889 ? (((a ? a : 6522) | (a & 14'd1837)) << 2) : 15912));
            
            default: result_0949 = 14'd6638;
        endcase
    end

endmodule
        