
module simple_alu_0702(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0702
);

    always @(*) begin
        case(op)
            
            4'd0: result_0702 = (14'd1413 | (14'd11908 ^ (14'd8366 << 3)));
            
            4'd1: result_0702 = (~(((a << 3) ^ (a ^ (b ^ 14'd12967))) & (~(b & (a ^ 14'd2837)))));
            
            4'd2: result_0702 = (~((14'd5745 + ((b & a) + (b * 14'd11944))) ^ (~14'd12517)));
            
            4'd3: result_0702 = (a | (14'd8663 << 1));
            
            4'd4: result_0702 = (14'd9014 ^ ((((14'd10853 << 3) >> 1) << 3) | (((14'd9599 << 2) << 2) >> 1)));
            
            4'd5: result_0702 = ((b | ((a + (~a)) - ((14'd1495 + a) * 14'd9692))) >> 3);
            
            4'd6: result_0702 = (((((14'd7390 + 14'd4797) << 3) >> 1) & (14'd12159 & ((14'd15604 - a) >> 3))) & (14'd739 >> 3));
            
            4'd7: result_0702 = ((((a ? (a >> 2) : 6454) - ((14'd8121 ? 14'd13352 : 14270) - 14'd7973)) >> 3) * (a - (((14'd6589 >> 2) - (14'd11862 * a)) | (~14'd5519))));
            
            4'd8: result_0702 = (((~(~(a | 14'd5842))) >> 3) ? b : 6763);
            
            4'd9: result_0702 = (14'd8279 >> 3);
            
            4'd10: result_0702 = (~(((14'd7242 << 3) & ((a ? 14'd6032 : 15870) + (~a))) * ((14'd1281 * (14'd5588 * 14'd11830)) >> 3)));
            
            4'd11: result_0702 = (14'd2823 | (14'd6831 << 3));
            
            4'd12: result_0702 = ((b * (b & ((14'd10295 + 14'd2788) | b))) | ((((14'd7150 ^ a) ^ (~14'd1533)) & ((b ^ b) ^ 14'd4676)) * (((14'd2677 - a) ^ b) + (a & (b + 14'd4553)))));
            
            default: result_0702 = a;
        endcase
    end

endmodule
        