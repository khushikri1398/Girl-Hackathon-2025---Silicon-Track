
module simple_alu_0138(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0138
);

    always @(*) begin
        case(op)
            
            4'd0: result_0138 = (((((14'd7113 & 14'd2367) - (14'd4690 & 14'd2370)) + ((~a) + (14'd12477 - a))) >> 2) << 2);
            
            4'd1: result_0138 = (a ^ (b | (((14'd9294 >> 2) + (~b)) & b)));
            
            4'd2: result_0138 = (~14'd10138);
            
            4'd3: result_0138 = (~(((a - (14'd11456 & 14'd14651)) << 3) ^ (((14'd8421 >> 3) ^ (14'd1746 + b)) ^ ((14'd5488 << 2) << 1))));
            
            4'd4: result_0138 = (((~((14'd737 ^ 14'd254) & b)) << 1) >> 3);
            
            4'd5: result_0138 = ((((b >> 2) + ((14'd7888 - b) & b)) - ((14'd16156 * (~b)) ? ((14'd2239 ? a : 1217) | a) : 14335)) * 14'd8130);
            
            4'd6: result_0138 = (((a | ((a * a) + (a & 14'd16329))) + 14'd3327) | (~((14'd6668 >> 1) >> 1)));
            
            default: result_0138 = 14'd415;
        endcase
    end

endmodule
        