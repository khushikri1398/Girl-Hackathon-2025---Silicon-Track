
module simple_alu_0637(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0637
);

    always @(*) begin
        case(op)
            
            4'd0: result_0637 = (a + ((((14'd4494 >> 3) >> 3) - ((14'd2702 - b) | (14'd3273 * 14'd3265))) | (((a ? 14'd9464 : 142) ^ (14'd2331 & 14'd10427)) << 3)));
            
            4'd1: result_0637 = (((a | (~(~14'd969))) << 1) | ((((14'd11615 ^ 14'd2081) - (14'd13162 & 14'd5106)) + (~(14'd16158 & 14'd11567))) >> 1));
            
            4'd2: result_0637 = (((((~b) ^ (14'd8927 ? b : 5009)) ^ ((~a) << 1)) << 3) >> 2);
            
            4'd3: result_0637 = (((((14'd4887 | b) + b) - ((14'd2264 >> 3) - (a ^ 14'd7215))) + (((~14'd14311) + (14'd10617 * b)) << 3)) & (((a ^ (14'd6773 * 14'd11726)) ? (b & (b * 14'd10833)) : 917) - (~14'd2971)));
            
            4'd4: result_0637 = ((14'd4753 | 14'd2545) * b);
            
            4'd5: result_0637 = (14'd13708 - (14'd14983 << 1));
            
            4'd6: result_0637 = (((((~b) + a) ^ ((14'd7872 ? b : 9260) >> 1)) + (((b ^ 14'd12013) | (14'd11419 ? 14'd9928 : 9272)) & 14'd16274)) | (((a ^ (b << 3)) >> 3) * (~(~(a ? 14'd10690 : 11367)))));
            
            4'd7: result_0637 = (~(((14'd13060 ? (14'd416 >> 1) : 11524) | (14'd4629 + (b + 14'd13745))) << 2));
            
            4'd8: result_0637 = (14'd7473 << 2);
            
            4'd9: result_0637 = (~b);
            
            4'd10: result_0637 = (~((~(b + (14'd13196 & b))) ? 14'd12657 : 11564));
            
            4'd11: result_0637 = (((~14'd14542) ? ((~(b + b)) << 2) : 12229) >> 2);
            
            4'd12: result_0637 = ((b ? 14'd15837 : 15552) & b);
            
            4'd13: result_0637 = (14'd2564 << 3);
            
            4'd14: result_0637 = (((14'd2443 ^ ((14'd16114 ? 14'd11786 : 7238) << 2)) * (14'd14545 + 14'd4797)) ? ((~((b * b) | (14'd2978 >> 2))) | (a ? (14'd14665 * (b ^ b)) : 643)) : 6298);
            
            default: result_0637 = 14'd1785;
        endcase
    end

endmodule
        