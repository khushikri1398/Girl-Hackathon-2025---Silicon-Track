
module simple_alu_0037(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0037
);

    always @(*) begin
        case(op)
            
            4'd0: result_0037 = (b - 14'd14518);
            
            4'd1: result_0037 = ((~(((~a) << 2) & 14'd15593)) ? ((a & (~(14'd4409 | 14'd14457))) - (((14'd7511 * 14'd14666) << 2) - ((b + 14'd3734) ? b : 12300))) : 4982);
            
            4'd2: result_0037 = (14'd7065 ? b : 14012);
            
            4'd3: result_0037 = ((((~(14'd5620 ^ b)) * 14'd12666) - 14'd3967) >> 3);
            
            4'd4: result_0037 = ((((~14'd7957) | 14'd10376) - 14'd13223) - (b | 14'd217));
            
            4'd5: result_0037 = (~((a - ((~14'd4500) + (14'd5124 + 14'd9154))) + (((b ^ b) & (14'd4605 ? b : 11395)) & 14'd942)));
            
            4'd6: result_0037 = ((a ^ 14'd4902) >> 2);
            
            4'd7: result_0037 = (((((14'd7455 + b) >> 1) << 2) & ((~14'd2199) >> 3)) * (~a));
            
            4'd8: result_0037 = (a - ((((14'd4963 >> 2) - (14'd4412 << 1)) << 2) - 14'd14669));
            
            4'd9: result_0037 = (~a);
            
            4'd10: result_0037 = (((((~14'd14094) ^ (a >> 2)) - ((14'd9872 >> 1) ? (14'd4943 * 14'd12118) : 3053)) | ((a * (14'd13632 ^ a)) | ((b + 14'd12191) * (a + 14'd14476)))) - (((~(~b)) | ((14'd7581 << 3) * (14'd14430 | 14'd4222))) * (((14'd3106 & b) * (14'd6104 >> 2)) | ((14'd6804 >> 3) & (a & b)))));
            
            default: result_0037 = b;
        endcase
    end

endmodule
        