
module simple_alu_0655(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0655
);

    always @(*) begin
        case(op)
            
            4'd0: result_0655 = (((((14'd6020 ? b : 6240) ? (14'd3621 ? 14'd2737 : 8366) : 3681) >> 2) ? ((~(14'd7643 | a)) - (~b)) : 15329) << 2);
            
            4'd1: result_0655 = (~((((14'd4632 | 14'd9096) + (~a)) << 2) & (a - ((a ? 14'd1337 : 9070) << 2))));
            
            4'd2: result_0655 = ((((b << 3) << 3) | (14'd15097 << 3)) * 14'd9367);
            
            4'd3: result_0655 = (((((14'd8199 * b) ? (14'd2468 ? 14'd3809 : 15912) : 11043) + ((14'd12222 >> 1) - (14'd5151 ^ 14'd14429))) + ((~14'd2590) + ((14'd12468 & 14'd5732) | (~a)))) << 3);
            
            4'd4: result_0655 = (((14'd9159 << 3) ? ((14'd8869 - b) ^ ((14'd14049 ? 14'd1223 : 999) | (a ^ 14'd8194))) : 3792) << 1);
            
            4'd5: result_0655 = (b + (((14'd9881 - (14'd5005 - 14'd4252)) + ((14'd13028 ^ 14'd9885) - b)) & ((b * 14'd14235) - ((b - 14'd11950) >> 3))));
            
            4'd6: result_0655 = ((~b) | ((((~14'd8465) | 14'd7240) & ((a << 3) | (14'd1935 ? b : 15425))) ^ a));
            
            4'd7: result_0655 = ((14'd4757 + (b | ((a ^ a) >> 1))) >> 2);
            
            4'd8: result_0655 = ((14'd1803 & (((~14'd5035) * (14'd11607 * 14'd2075)) * 14'd14340)) ? 14'd1272 : 4114);
            
            4'd9: result_0655 = ((14'd9072 ^ ((14'd6800 ^ 14'd3386) ^ ((14'd15739 | b) & (a << 2)))) - (14'd799 & 14'd16069));
            
            4'd10: result_0655 = (a >> 2);
            
            4'd11: result_0655 = (((~14'd15780) << 2) * 14'd3891);
            
            4'd12: result_0655 = ((~14'd15850) & ((((14'd5674 ^ 14'd13096) ^ (14'd1783 ? a : 2653)) * 14'd1092) ? (((a - 14'd15659) ? (b ^ 14'd7042) : 3386) * (a - (a >> 2))) : 15825));
            
            4'd13: result_0655 = ((14'd12561 << 1) | (14'd13082 + b));
            
            4'd14: result_0655 = (((~14'd1333) * (((14'd8705 >> 1) * (14'd3725 * 14'd11838)) + 14'd12656)) >> 3);
            
            default: result_0655 = a;
        endcase
    end

endmodule
        