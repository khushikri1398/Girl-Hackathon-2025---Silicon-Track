
module simple_alu_0991(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0991
);

    always @(*) begin
        case(op)
            
            4'd0: result_0991 = ((((a ^ (14'd8338 & b)) ^ ((14'd598 - 14'd1191) * 14'd6529)) * (((14'd2684 ^ 14'd4660) - (a | 14'd5501)) ? (~a) : 9266)) + (((14'd3733 & (14'd11899 & 14'd11841)) | ((14'd3960 & a) >> 2)) >> 2));
            
            4'd1: result_0991 = ((~(((14'd13241 ? b : 13750) + (a * a)) ^ ((14'd6090 * 14'd6784) ^ (b * 14'd314)))) & (((a << 3) >> 2) ^ 14'd3943));
            
            4'd2: result_0991 = ((b - 14'd6399) << 3);
            
            4'd3: result_0991 = ((a << 3) & 14'd16045);
            
            4'd4: result_0991 = (((14'd1819 - ((a >> 1) + (14'd957 | 14'd6073))) >> 3) ^ ((((14'd13473 ? 14'd820 : 10004) | (14'd9467 ? 14'd3702 : 3976)) - ((14'd9298 & b) | (a + a))) << 1));
            
            4'd5: result_0991 = (14'd8831 << 1);
            
            4'd6: result_0991 = (((((a | 14'd11379) - 14'd1119) ? ((14'd13566 << 3) ? b : 884) : 7497) >> 2) * (~a));
            
            4'd7: result_0991 = ((~(((14'd9426 << 1) >> 1) & ((14'd5365 & a) | b))) + (((a << 1) - ((14'd11725 - 14'd2638) - (a ? a : 15262))) << 3));
            
            4'd8: result_0991 = (~14'd4312);
            
            4'd9: result_0991 = (14'd11933 | ((~(a | a)) << 2));
            
            4'd10: result_0991 = (((~(~(14'd4289 >> 3))) << 1) * a);
            
            4'd11: result_0991 = (14'd3761 * ((((b & b) << 3) * ((a ? b : 13167) - (14'd779 | 14'd13088))) * ((~(a << 3)) - ((14'd10963 << 1) + a))));
            
            4'd12: result_0991 = (a | a);
            
            4'd13: result_0991 = (14'd11753 >> 2);
            
            4'd14: result_0991 = (14'd4234 - (~(b & (a | b))));
            
            4'd15: result_0991 = (((((b * 14'd9522) ^ (~14'd7915)) * (b >> 1)) | ((14'd2501 + (14'd15054 - b)) - (b * (14'd8315 >> 3)))) & a);
            
            default: result_0991 = 14'd14652;
        endcase
    end

endmodule
        