
module simple_alu_0486(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0486
);

    always @(*) begin
        case(op)
            
            4'd0: result_0486 = ((14'd7403 - 14'd12617) & 14'd12181);
            
            4'd1: result_0486 = (b ^ 14'd15281);
            
            4'd2: result_0486 = ((14'd15928 & 14'd884) + (((14'd13309 * (14'd2903 ? a : 15652)) | ((14'd3594 & b) + 14'd11249)) >> 3));
            
            4'd3: result_0486 = ((a ^ (((~b) + (~14'd147)) + (a & (14'd5471 | b)))) << 1);
            
            4'd4: result_0486 = (14'd8891 | (~(14'd11817 << 3)));
            
            4'd5: result_0486 = (((((a | b) + (b + b)) & ((14'd2476 ^ 14'd927) ? (14'd14895 * b) : 14670)) | (((14'd6205 | b) >> 1) + ((14'd13573 + 14'd3100) + 14'd12859))) - (((14'd14552 << 2) >> 3) ? (a - ((b >> 3) - 14'd3832)) : 3363));
            
            4'd6: result_0486 = ((a | ((a << 2) & ((a ? b : 1886) | b))) + ((((14'd8618 & 14'd9) - (a - b)) >> 2) - (((b | 14'd1063) ^ (~14'd5600)) >> 1)));
            
            4'd7: result_0486 = (14'd2675 - ((14'd11447 & ((14'd3623 * 14'd9347) | (a ^ 14'd16327))) | ((14'd11945 ^ a) ? (~b) : 6801)));
            
            4'd8: result_0486 = (~((14'd13598 - ((b << 2) << 1)) * ((~(b ^ a)) >> 1)));
            
            4'd9: result_0486 = (a ? (a ^ (((a ^ 14'd5237) * (a - 14'd5264)) * ((b | 14'd7751) - a))) : 3167);
            
            default: result_0486 = 14'd10354;
        endcase
    end

endmodule
        