
module simple_alu_0555(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0555
);

    always @(*) begin
        case(op)
            
            4'd0: result_0555 = (((((~b) & 14'd15938) ? (14'd15131 >> 3) : 1107) - ((14'd3006 | (14'd8420 >> 2)) - (a + (b >> 1)))) | b);
            
            4'd1: result_0555 = ((14'd9758 ^ (((14'd5074 | b) ? (a * 14'd14202) : 9719) * ((b & 14'd11201) ? 14'd14880 : 5937))) | ((~((14'd4860 + a) << 3)) + (((a ? 14'd7170 : 7396) - (b - a)) - ((14'd11033 - 14'd16122) + (14'd16078 * a)))));
            
            4'd2: result_0555 = (14'd6044 ^ a);
            
            4'd3: result_0555 = (14'd14557 >> 1);
            
            4'd4: result_0555 = (((b & ((14'd12816 ^ 14'd15892) + (a * 14'd438))) ? ((14'd1455 - (b + 14'd6936)) << 1) : 12097) ? ((((14'd499 | b) >> 3) * ((14'd1253 & 14'd4752) << 2)) & ((14'd11104 >> 2) << 2)) : 12904);
            
            4'd5: result_0555 = (~((((14'd11338 << 2) ? 14'd4290 : 14447) * ((b + 14'd15093) | (14'd9955 ^ 14'd9339))) * (14'd5903 | ((b & b) | (~14'd12404)))));
            
            4'd6: result_0555 = (14'd15327 ? (((a - 14'd9362) ^ ((14'd11695 >> 1) >> 2)) ? (~((14'd14086 | b) + 14'd10146)) : 1495) : 2757);
            
            4'd7: result_0555 = (((14'd6504 ? ((14'd224 - b) ^ 14'd14438) : 13926) ? 14'd11901 : 11300) ^ ((b | ((14'd13951 ? a : 16035) >> 3)) ? (14'd11753 >> 3) : 980));
            
            4'd8: result_0555 = ((~((14'd3286 | 14'd6436) ? ((14'd11345 ? b : 10619) << 3) : 2533)) - ((((14'd14133 | 14'd3745) * a) >> 3) - (b >> 2)));
            
            4'd9: result_0555 = (a & (14'd6489 << 2));
            
            4'd10: result_0555 = (~(~(14'd3822 | ((14'd12096 >> 2) - (b >> 3)))));
            
            4'd11: result_0555 = ((14'd11543 ^ (((a << 2) >> 3) >> 1)) + 14'd5642);
            
            default: result_0555 = b;
        endcase
    end

endmodule
        