
module simple_alu_0764(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0764
);

    always @(*) begin
        case(op)
            
            4'd0: result_0764 = ((14'd10573 + (((~14'd14295) << 2) & ((14'd2318 + 14'd12749) ? (~14'd11018) : 3733))) & 14'd4000);
            
            4'd1: result_0764 = (((((14'd4411 + 14'd2116) << 1) << 1) ^ (b - ((b >> 2) * (a ? 14'd9274 : 4650)))) + (a * 14'd14075));
            
            4'd2: result_0764 = ((14'd7511 ^ (((b | 14'd14848) & (14'd10123 << 2)) >> 1)) ^ b);
            
            4'd3: result_0764 = (14'd1469 ^ b);
            
            4'd4: result_0764 = ((14'd11013 | ((14'd6534 + (a >> 1)) & ((14'd8561 & 14'd3687) << 3))) & b);
            
            4'd5: result_0764 = ((((14'd8373 - (b << 3)) & 14'd10914) + (((14'd10454 & a) - 14'd6731) | (a - 14'd1801))) + (a ^ 14'd4734));
            
            4'd6: result_0764 = (b | 14'd15299);
            
            default: result_0764 = 14'd15646;
        endcase
    end

endmodule
        