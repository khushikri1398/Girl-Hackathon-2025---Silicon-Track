
module simple_alu_0716(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0716
);

    always @(*) begin
        case(op)
            
            4'd0: result_0716 = ((b ^ (((14'd9795 >> 3) + (a << 2)) & 14'd5073)) * 14'd2089);
            
            4'd1: result_0716 = ((~((~(b << 3)) - 14'd356)) * (b * (~((b >> 1) + (b * 14'd3229)))));
            
            4'd2: result_0716 = (((14'd11586 ? ((14'd11421 - b) + 14'd6328) : 9494) & 14'd12927) | (a * 14'd7016));
            
            4'd3: result_0716 = (14'd3600 ? ((((14'd4582 << 2) | (14'd11099 + a)) ^ ((14'd919 + 14'd7020) >> 1)) - (((~b) << 3) >> 1)) : 12778);
            
            4'd4: result_0716 = ((b - 14'd14676) >> 1);
            
            4'd5: result_0716 = (((14'd10807 << 1) * 14'd14172) * (((14'd4363 | (b ^ 14'd7406)) >> 3) & 14'd1312));
            
            4'd6: result_0716 = (b | ((b + ((14'd3924 - 14'd4088) << 1)) ? (b + ((b * 14'd402) << 3)) : 11941));
            
            4'd7: result_0716 = (((14'd7076 >> 3) + 14'd5342) - ((((14'd8732 * a) & a) >> 1) & (((14'd7088 - 14'd14577) & (b >> 3)) ? a : 14148)));
            
            4'd8: result_0716 = ((14'd3786 >> 2) >> 3);
            
            4'd9: result_0716 = ((14'd13904 ^ (((14'd15406 ^ 14'd8916) & (14'd11021 * 14'd632)) + b)) * ((((14'd9197 * 14'd11787) ^ 14'd8510) ^ (b * (b ? 14'd799 : 5203))) * (((~14'd9541) ^ (14'd12399 << 3)) * ((~14'd1391) >> 3))));
            
            4'd10: result_0716 = ((14'd8191 << 3) + 14'd1815);
            
            4'd11: result_0716 = ((((14'd8661 * (14'd7701 - 14'd2795)) >> 2) << 2) ^ ((~a) ? 14'd7851 : 6391));
            
            default: result_0716 = 14'd12226;
        endcase
    end

endmodule
        