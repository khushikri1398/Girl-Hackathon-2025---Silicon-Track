
module simple_alu_0283(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0283
);

    always @(*) begin
        case(op)
            
            4'd0: result_0283 = ((b * (((14'd9144 ^ 14'd4027) | (14'd3690 * b)) & (14'd12665 & (a + 14'd11633)))) ? b : 4327);
            
            4'd1: result_0283 = (14'd4264 * b);
            
            4'd2: result_0283 = ((14'd8866 << 3) | (a + (((14'd1312 - b) * (14'd7943 ^ 14'd12209)) & ((~14'd3051) & a))));
            
            4'd3: result_0283 = (((~((14'd10514 << 1) & (b << 2))) - (~(b ? (14'd8314 * 14'd4802) : 930))) & ((((14'd7402 & 14'd3760) << 1) + b) ^ (((14'd3068 & a) << 2) >> 2)));
            
            4'd4: result_0283 = (((((14'd12796 ^ 14'd10876) * (b << 2)) - 14'd11677) | (~(~a))) ^ 14'd4825);
            
            4'd5: result_0283 = (~(~14'd9632));
            
            4'd6: result_0283 = (((((14'd7246 << 3) & (14'd315 ? 14'd12489 : 12434)) ? ((14'd10050 + b) + 14'd2374) : 15437) ^ (((b >> 3) | (14'd10268 - a)) ? (~14'd7600) : 10017)) << 3);
            
            4'd7: result_0283 = ((14'd14226 + (14'd142 * ((14'd8179 - b) - 14'd4203))) ? ((((a >> 3) | 14'd10610) + 14'd5395) ? a : 6069) : 4413);
            
            4'd8: result_0283 = (((((14'd1822 ^ 14'd7220) & (14'd5403 ? 14'd10373 : 10583)) + ((~14'd11986) ^ (a - b))) & (~((14'd13466 | 14'd6151) >> 1))) & b);
            
            4'd9: result_0283 = (((((14'd8324 ? b : 8888) * (b - 14'd14068)) - 14'd12736) - b) & ((((a | 14'd14260) ^ (14'd9335 >> 2)) ^ 14'd9365) ^ (~b)));
            
            4'd10: result_0283 = (14'd657 + 14'd9328);
            
            4'd11: result_0283 = ((~(((14'd5956 ? b : 10003) >> 2) ? ((~b) & (b * a)) : 12276)) & 14'd7243);
            
            4'd12: result_0283 = ((~(((14'd4601 * a) - (a << 2)) * ((14'd5253 >> 1) >> 3))) ? ((14'd9687 - 14'd223) + ((14'd1980 ^ 14'd1759) | ((14'd6618 & 14'd3569) - (~a)))) : 178);
            
            4'd13: result_0283 = ((~(((a << 1) | (14'd12420 + a)) + ((~14'd1195) ? (14'd4211 | 14'd3018) : 4249))) | 14'd12921);
            
            default: result_0283 = a;
        endcase
    end

endmodule
        