
module simple_alu_0162(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0162
);

    always @(*) begin
        case(op)
            
            4'd0: result_0162 = (((((14'd4880 & 14'd4310) ^ (14'd13582 ? 14'd10030 : 4378)) - a) ^ (((14'd1861 - b) + (b | 14'd8162)) & (~(14'd12753 - b)))) >> 3);
            
            4'd1: result_0162 = ((((~(b | b)) ? ((14'd9391 ^ 14'd1470) | (~14'd9738)) : 2720) - (((14'd10584 * 14'd11590) - 14'd12305) & 14'd8847)) - (14'd10985 & 14'd7992));
            
            4'd2: result_0162 = (14'd10249 << 2);
            
            4'd3: result_0162 = ((((14'd3148 | (14'd857 ? 14'd15132 : 15956)) & ((14'd7203 + a) ? 14'd5803 : 15846)) << 2) ? (((14'd746 * (14'd14515 >> 1)) << 2) - (((14'd8785 - 14'd15410) - (14'd11774 - 14'd15788)) ? (~(b + b)) : 10668)) : 2533);
            
            4'd4: result_0162 = (14'd15295 << 3);
            
            4'd5: result_0162 = ((14'd6532 ^ ((14'd9764 >> 3) - (~14'd15346))) - (((a << 1) ^ ((b ^ 14'd7293) * (14'd10193 ? 14'd4550 : 15648))) | (((14'd13604 << 2) ? (14'd2829 << 3) : 8337) * a)));
            
            4'd6: result_0162 = ((14'd814 | (b * ((b - a) & (a + 14'd16307)))) ? (~(((b | 14'd6811) * (14'd9228 ^ a)) >> 1)) : 6287);
            
            4'd7: result_0162 = (14'd700 ^ ((~((14'd8323 - 14'd541) & (14'd14436 >> 1))) << 3));
            
            4'd8: result_0162 = (b & (14'd11115 | (((a & b) >> 3) ? 14'd10328 : 523)));
            
            4'd9: result_0162 = (((b ^ 14'd6760) * (((14'd8437 - 14'd5663) & b) * (14'd11155 ^ (14'd5416 << 3)))) ^ (~((14'd6749 * (14'd6889 ? a : 46)) << 1)));
            
            4'd10: result_0162 = ((((a >> 2) | ((b * b) - (b >> 2))) | ((~14'd3131) >> 1)) | (14'd953 - (((b ^ 14'd6519) ^ (14'd5213 * a)) - 14'd480)));
            
            4'd11: result_0162 = (((a ^ 14'd3074) ^ ((14'd10381 ^ 14'd13174) | 14'd11946)) - ((14'd4264 & (a + (14'd4446 * 14'd6214))) ? (((b + a) - 14'd9210) << 2) : 6945));
            
            4'd12: result_0162 = ((~14'd4302) ? ((14'd9302 << 3) & 14'd13381) : 5434);
            
            4'd13: result_0162 = (~a);
            
            4'd14: result_0162 = (~(((14'd14639 & (14'd10672 << 1)) >> 1) ^ (((14'd12127 - 14'd12494) * (14'd8275 ^ b)) >> 1)));
            
            default: result_0162 = a;
        endcase
    end

endmodule
        