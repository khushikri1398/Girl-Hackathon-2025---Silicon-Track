
module simple_alu_0986(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0986
);

    always @(*) begin
        case(op)
            
            4'd0: result_0986 = (b & ((((14'd11556 << 1) << 1) | 14'd2663) | (((b + 14'd2930) - (14'd3856 | b)) ? a : 6734)));
            
            4'd1: result_0986 = (b * 14'd5909);
            
            4'd2: result_0986 = (((a ? (14'd7928 >> 2) : 795) >> 3) - ((((b * b) - (14'd15777 + 14'd8582)) | (b >> 1)) - (~((14'd15432 ? 14'd14373 : 5254) << 1))));
            
            4'd3: result_0986 = (((((a + 14'd6141) ? (b * 14'd10102) : 5156) ? (b & 14'd10415) : 73) | 14'd12497) << 2);
            
            4'd4: result_0986 = (((((14'd5708 ^ 14'd9551) << 1) | ((14'd15561 & 14'd16365) | a)) ? b : 345) - 14'd11173);
            
            4'd5: result_0986 = (~((~((b ? 14'd9401 : 1793) - (14'd864 + b))) >> 3));
            
            4'd6: result_0986 = ((14'd7120 << 3) * ((~((14'd16186 ^ 14'd2429) >> 2)) - 14'd2268));
            
            4'd7: result_0986 = ((~(((14'd16023 | 14'd8093) ? (14'd12496 ? 14'd11184 : 15021) : 5076) << 1)) ^ 14'd1449);
            
            4'd8: result_0986 = ((14'd8540 ? (((14'd9121 - 14'd7681) * a) << 2) : 14082) ^ 14'd3802);
            
            default: result_0986 = 14'd14677;
        endcase
    end

endmodule
        