
module simple_alu_0030(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0030
);

    always @(*) begin
        case(op)
            
            4'd0: result_0030 = (b + (a << 2));
            
            4'd1: result_0030 = ((((b - 12'd3444) - 12'd1835) * b) * (((12'd2390 ? 12'd322 : 824) >> 2) << 1));
            
            4'd2: result_0030 = ((~12'd617) & (a ^ ((b ^ 12'd1884) | (a + 12'd1202))));
            
            4'd3: result_0030 = ((((b - 12'd1702) ? b : 2985) << 3) >> 2);
            
            4'd4: result_0030 = (((a * (a << 2)) * 12'd3530) & (((a ? 12'd1061 : 170) - (~b)) << 1));
            
            4'd5: result_0030 = ((((~12'd840) + (b | 12'd1606)) + (12'd608 - (a * 12'd3996))) << 3);
            
            4'd6: result_0030 = ((((b | 12'd142) * (~12'd1479)) >> 1) << 2);
            
            4'd7: result_0030 = (12'd3783 >> 2);
            
            4'd8: result_0030 = ((((a & a) | 12'd1075) * b) | a);
            
            4'd9: result_0030 = (a & ((12'd871 - (b ^ 12'd1677)) << 1));
            
            4'd10: result_0030 = (~12'd2503);
            
            4'd11: result_0030 = ((((12'd1170 >> 1) - (12'd2148 ^ 12'd2693)) * 12'd1879) * (((12'd2449 + 12'd2765) ^ a) * ((12'd166 * 12'd494) << 2)));
            
            4'd12: result_0030 = (b - 12'd2831);
            
            4'd13: result_0030 = (~(((12'd306 << 1) ? 12'd564 : 2988) ^ 12'd780));
            
            default: result_0030 = a;
        endcase
    end

endmodule
        