
module simple_alu_0040(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0040
);

    always @(*) begin
        case(op)
            
            4'd0: result_0040 = (((((14'd7279 + b) - 14'd972) | ((14'd10336 & 14'd4494) * (14'd2480 * b))) + a) & 14'd2328);
            
            4'd1: result_0040 = (((14'd627 ? ((14'd7919 ^ 14'd8576) + (14'd4575 ? 14'd6358 : 16279)) : 6132) | 14'd3089) ? a : 14053);
            
            4'd2: result_0040 = (((14'd6550 * ((14'd5972 | 14'd5754) | (14'd15465 + a))) ? b : 15982) + ((((14'd9776 * b) ? (14'd10071 >> 1) : 8596) + 14'd8822) + (b ? ((a >> 3) << 1) : 791)));
            
            4'd3: result_0040 = (((((14'd12912 - b) | (~14'd1426)) | (14'd6957 ? 14'd16356 : 8005)) >> 1) + (((14'd2431 + (14'd7053 - a)) << 2) * (~((14'd12910 & 14'd9107) | (b | 14'd14552)))));
            
            4'd4: result_0040 = (a ^ 14'd5242);
            
            4'd5: result_0040 = ((((14'd2876 ^ (14'd4983 | 14'd8416)) - ((14'd16171 ? a : 15314) ? 14'd362 : 3259)) ? (((~a) ^ (14'd13130 ? 14'd4197 : 4304)) ^ ((a * a) >> 1)) : 12980) >> 2);
            
            4'd6: result_0040 = ((((b * 14'd15844) & a) - b) ? (14'd9434 ^ (((14'd13498 * 14'd14372) + b) << 1)) : 12205);
            
            4'd7: result_0040 = (~((a ^ (~14'd2915)) * ((~14'd15986) | ((14'd3292 + a) >> 3))));
            
            4'd8: result_0040 = (((((a & 14'd16139) ^ (a * a)) & (b ^ (b << 1))) - a) - (14'd8050 ^ ((a ^ (14'd3810 & a)) | (14'd13723 | 14'd2852))));
            
            4'd9: result_0040 = (a ? ((14'd10770 << 3) + (((14'd15207 + 14'd11816) << 3) >> 3)) : 16245);
            
            default: result_0040 = 14'd1185;
        endcase
    end

endmodule
        