
module simple_alu_0251(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0251
);

    always @(*) begin
        case(op)
            
            4'd0: result_0251 = (b + (b | ((12'd1180 - a) & (b + 12'd428))));
            
            4'd1: result_0251 = (((12'd2136 << 2) * (b >> 3)) & (((12'd708 ^ b) + (a ^ 12'd3697)) & (12'd3331 << 2)));
            
            4'd2: result_0251 = ((((12'd1325 * b) ? (12'd810 >> 3) : 2761) ? ((~12'd997) & (12'd4061 & a)) : 163) * ((12'd1967 ? (~b) : 1813) * 12'd2945));
            
            4'd3: result_0251 = ((((~12'd353) | (~a)) ? ((b - 12'd3545) ^ (12'd2400 * b)) : 2353) ^ (~a));
            
            4'd4: result_0251 = ((((12'd1188 - b) | (12'd4055 + 12'd89)) ? b : 2739) | ((b << 2) + b));
            
            4'd5: result_0251 = ((12'd562 + (12'd455 | 12'd1874)) >> 1);
            
            4'd6: result_0251 = (((~(b - 12'd153)) * (~(b | a))) * a);
            
            4'd7: result_0251 = ((~a) + (((12'd1690 | 12'd2387) ? (b << 2) : 28) * ((12'd2869 - 12'd3458) | 12'd1446)));
            
            4'd8: result_0251 = ((12'd1896 ? ((~12'd2324) - 12'd1393) : 1352) >> 2);
            
            4'd9: result_0251 = ((((12'd906 << 3) & (12'd2561 ^ 12'd2552)) * (12'd3268 ^ (b ? 12'd1386 : 300))) >> 3);
            
            4'd10: result_0251 = (((~(12'd3584 - 12'd2323)) ? ((12'd1167 ? a : 1577) * (b << 1)) : 942) & (((b ? b : 1180) ? (12'd3991 * a) : 1368) - (12'd3936 >> 1)));
            
            4'd11: result_0251 = ((12'd3158 ^ ((12'd3327 ? b : 1326) | (b ^ a))) & 12'd3258);
            
            default: result_0251 = b;
        endcase
    end

endmodule
        