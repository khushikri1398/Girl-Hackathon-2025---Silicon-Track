
module simple_alu_0897(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0897
);

    always @(*) begin
        case(op)
            
            4'd0: result_0897 = (b - (b ? (14'd13450 >> 2) : 8970));
            
            4'd1: result_0897 = ((~a) ^ ((~(14'd8668 << 2)) | (((a + 14'd15375) - (14'd9175 - b)) ? ((b | 14'd13422) ? (14'd8843 | b) : 7859) : 9583)));
            
            4'd2: result_0897 = (~(~(14'd2211 & (14'd12906 << 2))));
            
            4'd3: result_0897 = (((a - ((14'd6966 - 14'd7982) + (~b))) * (14'd2052 ? ((14'd4149 << 2) ^ (~14'd6398)) : 10823)) * (14'd7815 ^ (14'd16264 & 14'd4322)));
            
            4'd4: result_0897 = ((14'd10207 >> 3) * b);
            
            4'd5: result_0897 = ((14'd7729 + ((~(b ^ b)) << 3)) & (((~(14'd11733 ^ 14'd1263)) * ((14'd6164 ? 14'd13123 : 6791) ^ (14'd7545 - 14'd12579))) & (((a - 14'd15443) - (14'd11549 >> 1)) - (b | (b * b)))));
            
            4'd6: result_0897 = (((((a + 14'd14339) >> 3) & (~(14'd6098 >> 2))) ^ ((~(14'd444 ? a : 3570)) ? (14'd2063 >> 1) : 14370)) & (a & (14'd6692 | a)));
            
            4'd7: result_0897 = (14'd2716 - (((14'd3077 ^ (b ^ a)) << 2) & (b + (a & (a ^ b)))));
            
            4'd8: result_0897 = (((((a >> 3) + (~b)) ? ((14'd5885 - 14'd1811) | (~14'd13032)) : 476) >> 1) | (((14'd4911 ? (14'd4976 | 14'd3823) : 1729) * ((14'd16034 >> 1) << 1)) ? (~((14'd8624 ? 14'd272 : 12968) ^ (~b))) : 14002));
            
            4'd9: result_0897 = (((((14'd4955 | 14'd11597) & (14'd7076 | b)) + a) - (((14'd834 ^ 14'd11147) | (~a)) + 14'd11814)) << 3);
            
            default: result_0897 = 14'd1285;
        endcase
    end

endmodule
        