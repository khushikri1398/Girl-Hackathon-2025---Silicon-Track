
module simple_alu_0966(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0966
);

    always @(*) begin
        case(op)
            
            4'd0: result_0966 = ((((14'd11779 + (14'd10630 << 3)) - ((14'd10112 * 14'd15650) | (a & 14'd2572))) ^ a) * ((14'd5518 * ((14'd10126 ^ 14'd5117) ? (b >> 1) : 13598)) + (14'd15649 | ((14'd8647 + b) + a))));
            
            4'd1: result_0966 = (((b >> 2) ^ 14'd5461) ^ 14'd6078);
            
            4'd2: result_0966 = (((((14'd310 + 14'd2677) ^ (a << 3)) - b) & (((14'd3784 - a) ^ (a ^ a)) + (~(a ^ 14'd4847)))) - ((((b * 14'd5022) >> 3) & 14'd4340) - (((14'd8747 * a) & (b - b)) * ((14'd3174 & 14'd15073) + (a + 14'd966)))));
            
            4'd3: result_0966 = ((14'd5440 * (((14'd9003 << 1) ? (14'd15980 << 1) : 15929) + (~(~14'd5420)))) << 1);
            
            4'd4: result_0966 = (14'd3703 >> 1);
            
            4'd5: result_0966 = (((b ? ((b ? 14'd10159 : 13561) + 14'd12944) : 14369) + (((14'd1348 + 14'd11981) >> 3) + 14'd461)) ? 14'd14864 : 7537);
            
            4'd6: result_0966 = (a >> 3);
            
            4'd7: result_0966 = (14'd2289 >> 2);
            
            4'd8: result_0966 = ((((a + a) >> 1) - 14'd11848) >> 1);
            
            4'd9: result_0966 = ((((a - (14'd1536 ^ 14'd12456)) ^ ((a << 3) | (14'd5873 ^ b))) ^ (((~a) >> 3) - (~(14'd1193 >> 1)))) ? (((b & 14'd11793) ? ((b & b) & (b >> 1)) : 4493) >> 3) : 10851);
            
            4'd10: result_0966 = (b - (((14'd1363 << 3) ? (14'd5965 & b) : 10066) * (14'd8491 ? ((14'd163 << 3) << 2) : 5846)));
            
            4'd11: result_0966 = (~((((a & 14'd13355) * (a * 14'd418)) ? ((b >> 1) ^ (a ^ 14'd14390)) : 15373) ? (~((14'd5887 | 14'd781) & (14'd4767 ^ b))) : 12415));
            
            4'd12: result_0966 = (((~((14'd6117 ? 14'd4608 : 10006) ? a : 8528)) | 14'd12322) >> 3);
            
            4'd13: result_0966 = (~((~14'd3356) ^ (((14'd7887 + 14'd11394) << 3) - (14'd272 >> 1))));
            
            default: result_0966 = 14'd12075;
        endcase
    end

endmodule
        