
module simple_alu_0936(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0936
);

    always @(*) begin
        case(op)
            
            4'd0: result_0936 = ((((~(b & 14'd1946)) - ((~a) ^ 14'd11703)) * ((14'd4071 & (14'd6916 ^ 14'd11192)) - (14'd12497 | (~a)))) * (((~(14'd4520 >> 3)) << 3) + a));
            
            4'd1: result_0936 = (~(~(((14'd3916 * a) >> 2) & ((14'd16113 - 14'd933) - (14'd6467 << 1)))));
            
            4'd2: result_0936 = (((14'd2047 + (~(a ? 14'd12104 : 8411))) | a) ^ (14'd13551 & 14'd6054));
            
            4'd3: result_0936 = ((~14'd6502) << 2);
            
            4'd4: result_0936 = ((14'd3126 ? 14'd12627 : 9687) ? ((((14'd7548 & 14'd15507) + (14'd14889 + 14'd5047)) ^ ((~14'd2416) >> 2)) + (~((b + 14'd13564) ? (14'd12534 ^ b) : 1081))) : 956);
            
            4'd5: result_0936 = (b ^ ((14'd2364 | (~(14'd5710 << 1))) >> 3));
            
            4'd6: result_0936 = (((14'd9973 - (b + 14'd0)) >> 1) << 1);
            
            4'd7: result_0936 = (((~a) | ((14'd4590 & (14'd1004 ^ 14'd4077)) ? (14'd10510 ? (a ? a : 11440) : 15444) : 15804)) ? (~(((14'd4620 & a) + (14'd383 & a)) & (a >> 3))) : 7636);
            
            4'd8: result_0936 = (14'd3561 ? (14'd2132 ? (((14'd13824 << 1) >> 3) ? (~(b ? 14'd5187 : 6757)) : 8758) : 8377) : 15682);
            
            4'd9: result_0936 = (~a);
            
            4'd10: result_0936 = ((14'd13594 | (14'd14142 | ((14'd7941 + 14'd13191) | (14'd11833 | a)))) * ((14'd907 ^ ((14'd14543 & a) << 2)) << 1));
            
            4'd11: result_0936 = (a & (14'd5369 - (((a & b) ? (b - b) : 2219) << 3)));
            
            4'd12: result_0936 = (~14'd1507);
            
            4'd13: result_0936 = (((((14'd10096 << 2) - (b << 3)) & (~(14'd8427 | a))) - a) ? ((((a * b) << 2) & ((a >> 2) + (14'd2055 * b))) - (((~b) ^ (14'd3084 * 14'd12066)) | b)) : 9864);
            
            4'd14: result_0936 = ((14'd13246 + (((14'd6470 + 14'd245) * (b ^ a)) | ((14'd3603 >> 2) >> 3))) | a);
            
            4'd15: result_0936 = ((14'd10109 | (((a + 14'd6102) | (14'd15387 | 14'd2607)) >> 2)) ^ (a + 14'd15264));
            
            default: result_0936 = 14'd7138;
        endcase
    end

endmodule
        