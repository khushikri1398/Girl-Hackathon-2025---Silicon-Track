
module simple_alu_0438(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0438
);

    always @(*) begin
        case(op)
            
            4'd0: result_0438 = ((b & a) ? b : 6242);
            
            4'd1: result_0438 = ((14'd3307 + (a + ((14'd15039 - 14'd2832) << 2))) + ((~(14'd12881 * (a ^ 14'd14505))) - ((b ? 14'd10241 : 11586) | (b >> 1))));
            
            4'd2: result_0438 = (((~((~14'd4242) - (14'd186 | b))) + ((14'd6297 >> 1) << 2)) - 14'd6223);
            
            4'd3: result_0438 = (((((14'd4793 | b) << 2) & (14'd12050 ? (b | a) : 1220)) * (((a * 14'd7929) * 14'd14374) | (~b))) - a);
            
            4'd4: result_0438 = (a * (~14'd7186));
            
            4'd5: result_0438 = (14'd9327 * ((((b & b) & (14'd853 & a)) ^ (b & (14'd973 - 14'd8116))) * (((14'd1832 ? 14'd13512 : 11266) + b) | (14'd119 | (14'd5255 + 14'd1992)))));
            
            4'd6: result_0438 = (((((b << 1) - (b - 14'd11343)) ? ((14'd15887 & a) | (14'd7361 << 2)) : 3415) & (~((~14'd5157) << 3))) ? ((((b & 14'd10080) * (14'd8515 * 14'd10136)) & ((14'd11873 & 14'd1465) & (14'd12859 ? a : 2497))) << 1) : 479);
            
            4'd7: result_0438 = (a + (~(((~b) + (14'd14515 ^ 14'd1160)) * ((14'd65 ? b : 1658) | (a >> 3)))));
            
            4'd8: result_0438 = ((14'd4632 << 1) - a);
            
            4'd9: result_0438 = ((14'd1531 * (a << 3)) + 14'd16057);
            
            4'd10: result_0438 = (((((14'd13265 | b) << 1) ? ((14'd12886 >> 1) << 2) : 9574) ? 14'd6699 : 10103) | ((((14'd12436 >> 1) & (b ? a : 8277)) - ((b ^ 14'd7810) ? (14'd579 + 14'd11319) : 4964)) + (~(b << 1))));
            
            default: result_0438 = 14'd9838;
        endcase
    end

endmodule
        