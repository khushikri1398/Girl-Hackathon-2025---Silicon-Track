
module simple_alu_0751(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0751
);

    always @(*) begin
        case(op)
            
            4'd0: result_0751 = ((((14'd13969 * 14'd12285) | ((14'd281 + 14'd391) + 14'd16111)) - (((a - a) << 1) ^ ((14'd1678 & b) << 2))) << 3);
            
            4'd1: result_0751 = (((((b - b) ^ (14'd1575 ^ a)) ? a : 6089) << 2) >> 3);
            
            4'd2: result_0751 = ((~(~((14'd6646 | b) >> 2))) | ((14'd5394 ? 14'd5362 : 1366) << 1));
            
            4'd3: result_0751 = (((a - b) ? (14'd2589 ^ ((14'd15719 - a) * 14'd3958)) : 1637) ? b : 13198);
            
            4'd4: result_0751 = (~14'd3885);
            
            4'd5: result_0751 = (~14'd11049);
            
            4'd6: result_0751 = ((~(((14'd2491 + a) * (~14'd823)) + (~(14'd9613 | 14'd15145)))) ^ ((14'd218 << 1) ^ (~((14'd9113 & 14'd2442) - (b + b)))));
            
            4'd7: result_0751 = ((b & (((14'd7195 * 14'd2266) + b) >> 2)) ? ((a ? ((14'd10928 - 14'd10061) + (a >> 1)) : 1501) - ((a | 14'd11594) << 3)) : 11730);
            
            4'd8: result_0751 = (((((14'd5844 ? a : 15587) ? (14'd2144 * 14'd7301) : 3805) * ((b - 14'd4398) ? (~14'd2543) : 4227)) & (((~14'd9070) >> 3) ? (14'd13223 << 2) : 4976)) + ((((b ? b : 9493) ? (14'd3876 >> 1) : 11747) >> 2) << 3));
            
            4'd9: result_0751 = ((14'd722 << 1) | ((((14'd2488 | 14'd7221) >> 2) >> 1) | (((~14'd13567) & (14'd12687 ? 14'd13347 : 12427)) * (~(14'd7568 ? a : 10488)))));
            
            4'd10: result_0751 = (((14'd12748 | (~(~14'd4255))) & (((14'd8111 - 14'd13745) ^ (14'd9022 ? 14'd1452 : 7201)) >> 2)) & (((14'd10594 << 1) * 14'd10283) + ((~(a & a)) + (14'd14894 & (14'd14841 * 14'd3044)))));
            
            4'd11: result_0751 = (14'd8556 >> 3);
            
            4'd12: result_0751 = (b & ((((14'd15996 * a) * (14'd12376 ^ 14'd2041)) << 1) ^ 14'd5247));
            
            default: result_0751 = 14'd849;
        endcase
    end

endmodule
        