
module simple_alu_0310(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0310
);

    always @(*) begin
        case(op)
            
            4'd0: result_0310 = (((~14'd843) + b) ? ((14'd7884 - 14'd4731) | b) : 10590);
            
            4'd1: result_0310 = ((14'd9213 ^ (((a - b) ? (14'd1650 - b) : 1947) << 2)) ^ (14'd8809 ? (14'd4266 ^ a) : 2575));
            
            4'd2: result_0310 = ((14'd10426 ? a : 16288) + ((((~a) | (14'd643 + 14'd10961)) & 14'd14524) + (((b | a) ^ (b ^ 14'd12939)) - ((14'd7270 & a) | 14'd7986))));
            
            4'd3: result_0310 = ((~(~14'd14087)) ? (a >> 1) : 7353);
            
            4'd4: result_0310 = ((14'd9337 + ((14'd2184 | (a | 14'd15091)) >> 2)) >> 3);
            
            4'd5: result_0310 = (((b ? (14'd12502 >> 3) : 1943) ? ((a & (14'd6261 >> 3)) | ((14'd9708 * b) * (14'd2485 ^ 14'd342))) : 14263) - (14'd2664 & (((14'd10667 ^ 14'd16333) >> 3) | 14'd10713)));
            
            4'd6: result_0310 = (((14'd7485 + 14'd12294) ? (((b | b) & 14'd10596) ^ (14'd2968 + (14'd8434 + b))) : 922) << 3);
            
            4'd7: result_0310 = (((~((a * 14'd4371) * b)) & 14'd8105) >> 3);
            
            4'd8: result_0310 = (~(14'd12484 >> 1));
            
            4'd9: result_0310 = (((((14'd10812 ? a : 2508) + 14'd14356) - ((14'd2017 - 14'd8916) << 3)) >> 3) >> 3);
            
            4'd10: result_0310 = (14'd11874 | (((14'd14148 & b) >> 2) | (14'd12444 + ((14'd4093 >> 3) ^ (14'd884 >> 2)))));
            
            4'd11: result_0310 = (a | b);
            
            4'd12: result_0310 = (((((14'd11436 | a) >> 1) | (14'd834 >> 1)) | ((14'd6313 * 14'd11673) | ((b >> 2) ^ (b >> 2)))) << 1);
            
            4'd13: result_0310 = ((~14'd8245) << 3);
            
            default: result_0310 = a;
        endcase
    end

endmodule
        