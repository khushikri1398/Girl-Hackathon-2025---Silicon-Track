
module simple_alu_0008(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0008
);

    always @(*) begin
        case(op)
            
            4'd0: result_0008 = ((~(a << 1)) >> 2);
            
            4'd1: result_0008 = ((14'd9525 ? 14'd8521 : 2311) ? ((((~14'd13694) >> 3) | ((14'd14770 << 1) ? (b ^ 14'd5698) : 8888)) >> 2) : 8928);
            
            4'd2: result_0008 = ((14'd12870 << 1) << 3);
            
            4'd3: result_0008 = (a ^ (((b * b) & (~(14'd14595 ^ 14'd11422))) << 2));
            
            4'd4: result_0008 = (((((14'd8162 ^ b) ? (14'd4583 << 2) : 9649) + 14'd14639) >> 2) & ((((b & b) ^ (14'd14919 | 14'd9058)) ^ 14'd6819) & ((~(14'd9564 ? 14'd5093 : 6310)) << 2)));
            
            4'd5: result_0008 = (((((~14'd11896) + (~14'd9732)) - (14'd4283 ^ 14'd12873)) << 2) ^ (14'd12091 * ((14'd3737 & (14'd5321 & 14'd14366)) ? a : 16100)));
            
            4'd6: result_0008 = (14'd15342 ? 14'd10674 : 8470);
            
            4'd7: result_0008 = (((((b << 2) - (14'd1105 & 14'd942)) + (14'd11191 | 14'd11020)) & 14'd691) - b);
            
            4'd8: result_0008 = (((((~a) >> 1) >> 2) & 14'd930) ? 14'd11730 : 3406);
            
            4'd9: result_0008 = (((((a - 14'd16231) + (14'd14075 ? 14'd8173 : 6533)) & (14'd5104 >> 1)) + (a | 14'd7164)) >> 2);
            
            default: result_0008 = 14'd10153;
        endcase
    end

endmodule
        