
module simple_alu_0711(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0711
);

    always @(*) begin
        case(op)
            
            4'd0: result_0711 = ((((14'd12726 >> 2) | ((14'd11127 ^ 14'd15868) ^ (a << 1))) >> 2) ^ (14'd8619 + (a & ((14'd11437 + b) + (b >> 2)))));
            
            4'd1: result_0711 = (((((a - b) ^ a) * 14'd8191) << 2) + 14'd11856);
            
            4'd2: result_0711 = (((~(b + (14'd14528 | b))) ^ 14'd9885) * ((14'd1234 * ((a + 14'd14394) >> 3)) * ((~14'd1995) + ((b | 14'd15931) >> 2))));
            
            4'd3: result_0711 = (((~((b | 14'd7015) - (14'd5598 + 14'd15346))) ^ (14'd6821 ^ ((14'd3037 << 3) - (14'd2140 ^ 14'd4535)))) | (((b & (14'd13836 & 14'd545)) ^ a) ? ((14'd8213 + (14'd2143 ^ 14'd6533)) + a) : 7474));
            
            4'd4: result_0711 = ((b >> 1) >> 1);
            
            4'd5: result_0711 = (14'd9732 ? ((~(14'd1866 + (14'd7060 >> 3))) * ((14'd13389 & a) ? (14'd5234 ? a : 7931) : 7779)) : 5401);
            
            4'd6: result_0711 = (((((14'd3236 | 14'd10940) * 14'd5727) >> 2) ^ 14'd11914) ? ((((b >> 3) * 14'd1163) ? ((~14'd12091) * (a >> 2)) : 6378) ^ 14'd7025) : 5448);
            
            4'd7: result_0711 = (((~b) << 3) & 14'd14324);
            
            4'd8: result_0711 = (~((((a << 3) | (14'd935 + 14'd7428)) ^ ((14'd8490 >> 2) + (14'd6423 ? 14'd3912 : 16158))) * b));
            
            4'd9: result_0711 = ((((b - 14'd772) << 2) << 1) - ((((14'd3584 - a) | (~14'd6674)) - ((14'd10898 ^ 14'd2047) ^ 14'd6501)) >> 1));
            
            4'd10: result_0711 = ((14'd8740 + (((b >> 1) ^ 14'd6016) | 14'd10041)) | ((14'd13940 & ((b + 14'd6747) - (14'd15619 | 14'd2464))) | (14'd10307 >> 3)));
            
            4'd11: result_0711 = (((14'd4653 << 3) * ((~(b * 14'd12774)) | 14'd3033)) - ((((~a) << 3) * (14'd12885 ? 14'd2257 : 15376)) << 1));
            
            default: result_0711 = a;
        endcase
    end

endmodule
        