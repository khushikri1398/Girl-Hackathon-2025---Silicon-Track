
module simple_alu_0537(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0537
);

    always @(*) begin
        case(op)
            
            4'd0: result_0537 = (((((~b) + (~14'd14009)) ? ((14'd2764 - a) ? (a ^ b) : 8301) : 5113) + 14'd15301) - (14'd16110 | (((a | 14'd12625) ? 14'd13166 : 14195) ^ ((14'd9146 << 3) & b))));
            
            4'd1: result_0537 = ((((b - (14'd15950 + 14'd12461)) * (a * (b << 1))) >> 1) - 14'd10570);
            
            4'd2: result_0537 = (14'd4524 ^ (14'd4490 - 14'd1405));
            
            4'd3: result_0537 = ((14'd4342 - (b - 14'd6322)) << 1);
            
            4'd4: result_0537 = (((((14'd14368 | 14'd1656) - (~a)) + ((14'd5374 * b) ^ (14'd12288 ^ 14'd14996))) ? (((14'd12359 ? 14'd5965 : 10944) >> 1) >> 3) : 2141) | a);
            
            4'd5: result_0537 = (((((b * a) * (a - 14'd11062)) | (~(14'd385 ? a : 1171))) - ((~b) << 3)) ? a : 12019);
            
            4'd6: result_0537 = (a + (14'd2344 & (14'd16293 >> 1)));
            
            4'd7: result_0537 = (a * (14'd10318 >> 1));
            
            4'd8: result_0537 = (b << 1);
            
            4'd9: result_0537 = (((~14'd1975) * (((14'd13750 & b) ^ (b >> 1)) & ((~14'd15012) >> 2))) & 14'd5379);
            
            4'd10: result_0537 = (b ^ 14'd5746);
            
            4'd11: result_0537 = (~b);
            
            4'd12: result_0537 = ((~(14'd16224 + (14'd5189 & b))) | (14'd1741 | (~(b + (a ^ 14'd3388)))));
            
            default: result_0537 = b;
        endcase
    end

endmodule
        