
module simple_alu_0372(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0372
);

    always @(*) begin
        case(op)
            
            4'd0: result_0372 = ((~14'd6119) | 14'd75);
            
            4'd1: result_0372 = (14'd7113 & (((14'd2812 & a) | ((14'd10258 + 14'd7234) & (14'd1506 * 14'd13694))) << 2));
            
            4'd2: result_0372 = (((((a | a) << 2) << 2) * 14'd3995) ? (~(a - (14'd7448 ^ (14'd8633 << 2)))) : 1558);
            
            4'd3: result_0372 = (((14'd13257 ^ (~(14'd8670 << 1))) * 14'd2057) - (~b));
            
            4'd4: result_0372 = (((a - a) * ((a ^ (14'd8900 << 2)) >> 1)) >> 1);
            
            4'd5: result_0372 = (((a >> 2) & ((b * (14'd9599 ^ 14'd13353)) ? 14'd10876 : 409)) & 14'd12707);
            
            default: result_0372 = b;
        endcase
    end

endmodule
        