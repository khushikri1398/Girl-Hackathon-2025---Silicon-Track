
module simple_alu_0476(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0476
);

    always @(*) begin
        case(op)
            
            4'd0: result_0476 = (14'd1815 + ((((14'd7613 - 14'd9660) | (a ? 14'd11262 : 7315)) - ((14'd8848 ^ 14'd11472) + (14'd9273 & 14'd12997))) ^ 14'd5359));
            
            4'd1: result_0476 = ((~14'd447) - (b >> 1));
            
            4'd2: result_0476 = ((14'd13133 - ((b - (b - a)) ^ ((~a) | (b >> 2)))) & (a | a));
            
            4'd3: result_0476 = ((14'd7931 << 2) + (14'd4445 >> 2));
            
            4'd4: result_0476 = (14'd13355 << 3);
            
            4'd5: result_0476 = ((a - ((14'd257 | (14'd7579 & 14'd10130)) << 3)) * (~(((a ^ 14'd663) ? (a >> 3) : 15493) ? ((14'd12800 ? 14'd10729 : 14274) << 2) : 4969)));
            
            4'd6: result_0476 = (14'd12177 * b);
            
            4'd7: result_0476 = ((~((14'd9819 ? b : 13429) ? ((~a) * (a >> 3)) : 10479)) + (((b - (b & a)) >> 1) ^ a));
            
            4'd8: result_0476 = ((14'd15191 * (14'd5617 >> 3)) << 1);
            
            4'd9: result_0476 = (14'd14853 - ((((14'd4024 | 14'd7950) * (14'd6660 ? a : 8076)) >> 1) - a));
            
            default: result_0476 = 14'd13478;
        endcase
    end

endmodule
        