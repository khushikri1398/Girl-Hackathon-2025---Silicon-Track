
module simple_alu_0014(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0014
);

    always @(*) begin
        case(op)
            
            4'd0: result_0014 = (~(14'd3529 ? (((~14'd12030) ^ (14'd13273 - 14'd2342)) * ((b << 2) << 1)) : 13698));
            
            4'd1: result_0014 = (~(((~(14'd4626 << 1)) ? (b ^ 14'd16062) : 6192) & 14'd7539));
            
            4'd2: result_0014 = (((((b ? 14'd1856 : 9865) << 2) | ((a - 14'd6761) ^ (b * 14'd6287))) + (((14'd2567 << 3) ^ (14'd8806 - 14'd1152)) ^ (14'd11189 - (b * 14'd14262)))) - (((~(14'd4961 | 14'd2122)) & (~a)) ? (14'd7664 << 1) : 7594));
            
            4'd3: result_0014 = ((((~(a ? 14'd408 : 15364)) >> 3) | ((~(14'd14467 ^ 14'd11727)) - (~(~14'd16014)))) | (((14'd7347 - (~14'd4616)) | 14'd11667) - (((14'd13213 | a) + 14'd110) + b)));
            
            4'd4: result_0014 = ((b - (((14'd6946 & b) ? (14'd9413 ? b : 11791) : 12141) >> 1)) | (a - (14'd1932 * ((14'd10492 & 14'd11723) >> 3))));
            
            4'd5: result_0014 = ((14'd1820 | (14'd15490 ^ ((~14'd10595) - a))) + 14'd11934);
            
            4'd6: result_0014 = ((a ? 14'd5759 : 1800) & 14'd16024);
            
            4'd7: result_0014 = (~((a + 14'd13718) - (((a ^ 14'd11241) + 14'd12452) ^ ((14'd13694 ^ a) << 1))));
            
            4'd8: result_0014 = (((((14'd3215 << 1) >> 3) + 14'd13777) >> 3) & (~(((14'd10897 ? 14'd874 : 4697) << 1) + (14'd10081 << 1))));
            
            4'd9: result_0014 = (a >> 2);
            
            4'd10: result_0014 = (14'd14198 + (14'd4909 | (((14'd11629 + 14'd7529) >> 1) ^ ((14'd13037 >> 2) & (~a)))));
            
            4'd11: result_0014 = (14'd6095 * (~(14'd10475 & (a << 2))));
            
            4'd12: result_0014 = (((((~14'd5502) ^ (b ? a : 7355)) & (a * (a + 14'd3446))) - 14'd6576) & (a + (14'd15236 >> 2)));
            
            4'd13: result_0014 = ((((14'd10740 ^ (a | 14'd7927)) >> 3) >> 1) ^ a);
            
            default: result_0014 = 14'd13199;
        endcase
    end

endmodule
        