
module simple_alu_0104(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0104
);

    always @(*) begin
        case(op)
            
            4'd0: result_0104 = ((a >> 1) ^ (14'd8099 >> 3));
            
            4'd1: result_0104 = (((14'd7090 | ((b ^ 14'd8021) ^ (~14'd7829))) << 1) - ((((14'd7336 - 14'd7281) >> 3) >> 3) & 14'd830));
            
            4'd2: result_0104 = ((((14'd920 + (14'd5939 * 14'd2170)) - (~b)) | (((~14'd869) >> 3) * ((~14'd14191) >> 1))) ^ 14'd11148);
            
            4'd3: result_0104 = (~((((14'd8487 ^ b) >> 1) - ((14'd7886 << 3) >> 3)) ^ 14'd14315));
            
            4'd4: result_0104 = ((a ^ (14'd13896 * ((14'd8145 * a) >> 3))) ? a : 1575);
            
            4'd5: result_0104 = (14'd4719 * ((((b - 14'd3143) + (b + a)) ? (a ? (14'd5423 ? b : 9427) : 4330) : 1005) + b));
            
            default: result_0104 = 14'd10580;
        endcase
    end

endmodule
        