
module simple_alu_0123(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0123
);

    always @(*) begin
        case(op)
            
            4'd0: result_0123 = (14'd12539 & (b >> 1));
            
            4'd1: result_0123 = (14'd4390 * (a - 14'd6313));
            
            4'd2: result_0123 = ((~(((~a) - (a << 3)) - 14'd26)) << 2);
            
            4'd3: result_0123 = (((14'd12384 * (14'd194 + (b | 14'd12879))) - (((14'd10561 >> 1) + 14'd221) ^ ((14'd2663 - 14'd5041) | (b >> 3)))) + 14'd12153);
            
            4'd4: result_0123 = ((((~(14'd8304 << 2)) * (a - 14'd8431)) ^ (a + ((14'd15227 * 14'd4465) | (b ? a : 7036)))) ? ((((14'd13886 | 14'd3302) - (14'd3957 ? a : 2578)) | ((14'd15886 + b) & b)) & (((14'd5599 ^ 14'd1820) - (b ^ b)) & ((14'd7593 ? 14'd14610 : 8798) - (14'd4037 << 3)))) : 3459);
            
            4'd5: result_0123 = (((((a + 14'd7073) >> 3) ^ ((14'd3783 & b) - (a >> 2))) * ((~(a | 14'd11771)) ^ (~(14'd3239 + a)))) | ((((~14'd4618) | (14'd2249 >> 1)) - ((14'd6493 | b) | 14'd13905)) & 14'd1539));
            
            4'd6: result_0123 = (b & ((((14'd4171 | 14'd11281) & 14'd766) ^ 14'd13601) | a));
            
            4'd7: result_0123 = (((((14'd1735 & 14'd7701) - 14'd575) * (14'd14229 * (14'd11951 >> 2))) ^ (14'd15280 - 14'd8931)) ? 14'd13684 : 11812);
            
            4'd8: result_0123 = (14'd7675 ^ (14'd15085 * 14'd5418));
            
            4'd9: result_0123 = ((14'd8915 >> 3) & (((14'd1989 & (b << 1)) ^ (14'd2618 ^ 14'd10095)) & ((~(~14'd6354)) << 2)));
            
            4'd10: result_0123 = ((~b) ? 14'd953 : 3965);
            
            4'd11: result_0123 = (14'd3906 << 3);
            
            4'd12: result_0123 = (((14'd1103 & ((14'd15421 + a) << 1)) ? (~(14'd6855 ^ b)) : 2949) + ((14'd4779 << 1) << 3));
            
            4'd13: result_0123 = (((14'd883 & 14'd4454) << 1) + b);
            
            4'd14: result_0123 = (((((14'd2549 + b) * (b | 14'd3261)) + (14'd12089 >> 2)) & a) ^ b);
            
            default: result_0123 = a;
        endcase
    end

endmodule
        