
module simple_alu_0375(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0375
);

    always @(*) begin
        case(op)
            
            4'd0: result_0375 = (((((b + b) + 14'd12807) - (14'd4571 - 14'd8361)) & (((a - 14'd1003) ^ a) - (~14'd788))) * ((b * ((a ^ 14'd10400) & 14'd11847)) >> 3));
            
            4'd1: result_0375 = ((((14'd2332 - (b >> 1)) ^ ((a * 14'd2406) >> 1)) + ((a << 1) + ((14'd14180 | a) >> 3))) ? (14'd8589 + a) : 3259);
            
            4'd2: result_0375 = (~((14'd3988 + ((14'd14294 + b) - (14'd1420 & 14'd8746))) | ((b | (b ^ 14'd10546)) ? ((b ^ b) ? (a << 3) : 4582) : 4606)));
            
            4'd3: result_0375 = ((~(((a + 14'd12774) + (b | 14'd13526)) - ((b >> 1) ^ a))) ? (~((14'd12479 ? (14'd8390 ? b : 6042) : 11483) | (14'd12192 ? (14'd3782 | 14'd11879) : 3458))) : 15652);
            
            default: result_0375 = a;
        endcase
    end

endmodule
        