
module simple_alu_0321(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0321
);

    always @(*) begin
        case(op)
            
            4'd0: result_0321 = ((14'd11708 + 14'd12687) - ((14'd3501 ^ (a | (14'd2878 + 14'd10684))) * 14'd1146));
            
            4'd1: result_0321 = (((~((14'd7127 * 14'd14881) & 14'd10331)) & 14'd13231) ^ (14'd2076 << 2));
            
            4'd2: result_0321 = (14'd8902 ? (a + (((b ? b : 10016) * (14'd6153 & 14'd10917)) * (14'd11017 << 2))) : 12261);
            
            4'd3: result_0321 = (b | 14'd7805);
            
            4'd4: result_0321 = (((((14'd4178 ^ b) >> 3) * ((~14'd4256) - (14'd8712 & b))) | a) << 3);
            
            4'd5: result_0321 = (((((14'd10075 >> 1) & (a + 14'd16044)) & ((a & a) << 3)) ? a : 10756) ? ((b - 14'd13666) + ((a - b) ? (b << 3) : 4651)) : 10853);
            
            4'd6: result_0321 = (14'd3264 - (((a ? (14'd2823 ? a : 15521) : 2363) << 2) - (((b - 14'd12501) & b) >> 1)));
            
            4'd7: result_0321 = (~b);
            
            4'd8: result_0321 = ((((14'd7022 << 3) << 3) ^ 14'd8993) ^ ((b & ((14'd9716 ^ b) * (14'd14105 << 2))) ^ (((14'd8978 << 1) ? (14'd1882 & a) : 6226) | 14'd2230)));
            
            4'd9: result_0321 = (((b << 3) ^ (((14'd6238 ^ 14'd11947) << 1) * ((a ? 14'd9110 : 12123) + 14'd5327))) - ((((b ^ b) ^ 14'd15281) | ((14'd926 + b) & b)) | (((14'd1738 * 14'd5025) * (~14'd7605)) >> 3)));
            
            4'd10: result_0321 = (~((((b + 14'd15403) + (a * 14'd14730)) ? (b | 14'd12046) : 1003) ? ((14'd13984 << 1) ? ((~14'd3151) ^ (14'd11713 - 14'd2592)) : 12270) : 13375));
            
            4'd11: result_0321 = (b << 1);
            
            4'd12: result_0321 = (14'd5869 ^ 14'd5782);
            
            4'd13: result_0321 = (((((14'd15185 + 14'd3241) * 14'd10189) * ((b * a) << 2)) ^ (14'd14007 * ((14'd7739 - 14'd8011) << 2))) * ((a >> 3) ^ ((14'd5757 | (14'd13250 | a)) | (14'd13135 * (~14'd10889)))));
            
            default: result_0321 = b;
        endcase
    end

endmodule
        