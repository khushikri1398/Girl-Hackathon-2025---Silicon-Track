
module simple_alu_0214(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0214
);

    always @(*) begin
        case(op)
            
            4'd0: result_0214 = ((b << 2) >> 2);
            
            4'd1: result_0214 = ((14'd11606 << 3) & ((((14'd4774 - b) >> 2) << 3) + a));
            
            4'd2: result_0214 = (((((~14'd11432) + 14'd15461) ^ (~(b ? 14'd5579 : 8405))) - ((~(a >> 3)) & ((14'd4881 + 14'd10361) * (14'd11395 ^ 14'd9904)))) & (~(((a ? b : 12078) << 1) | ((14'd9629 << 2) | (14'd8085 | 14'd1796)))));
            
            4'd3: result_0214 = (14'd1487 & 14'd363);
            
            4'd4: result_0214 = ((((14'd16249 << 2) << 1) + b) ^ ((((14'd4166 & 14'd9661) * (14'd16273 | a)) - a) ^ ((14'd6736 ^ (14'd5234 & a)) - ((a & a) >> 3))));
            
            4'd5: result_0214 = (b >> 3);
            
            default: result_0214 = 14'd1719;
        endcase
    end

endmodule
        