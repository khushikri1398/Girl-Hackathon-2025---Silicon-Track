
module simple_alu_0149(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0149
);

    always @(*) begin
        case(op)
            
            4'd0: result_0149 = ((((14'd13777 ? (14'd8617 - 14'd6742) : 7545) << 3) ^ (((14'd12278 ^ b) >> 3) + 14'd11438)) * ((14'd1489 - (~14'd14108)) + (14'd4238 ^ ((14'd14951 << 2) >> 1))));
            
            4'd1: result_0149 = (((((a * a) ^ (b * 14'd12890)) + ((~a) - (b ^ 14'd1138))) << 3) & (b * (~((14'd640 & 14'd11714) << 2))));
            
            4'd2: result_0149 = ((((~(14'd7950 & b)) | ((~14'd16212) >> 2)) * (((~b) ^ (b & a)) + ((b + 14'd12473) ? (14'd11416 >> 2) : 11193))) ^ (b & 14'd15644));
            
            4'd3: result_0149 = (14'd11126 - a);
            
            4'd4: result_0149 = ((14'd5489 ? a : 2451) + (((a + 14'd7814) << 3) | ((14'd16265 * (14'd9754 >> 1)) ? (14'd14919 + (14'd7658 - 14'd6488)) : 12786)));
            
            4'd5: result_0149 = ((a | (((a & 14'd479) - (14'd8539 + b)) | ((~14'd12442) + 14'd7591))) << 3);
            
            4'd6: result_0149 = (b * 14'd3837);
            
            4'd7: result_0149 = ((a * ((~(~b)) ? ((b * 14'd11420) - (14'd8259 ? 14'd7993 : 6151)) : 14017)) >> 3);
            
            4'd8: result_0149 = ((14'd477 * (b + 14'd12028)) ^ ((~((a >> 3) ^ (b ? 14'd2244 : 11469))) - (14'd1000 >> 1)));
            
            4'd9: result_0149 = (b ? (14'd11812 & 14'd2502) : 14209);
            
            4'd10: result_0149 = (a | 14'd648);
            
            4'd11: result_0149 = ((((a & 14'd9901) * ((a - b) | (14'd12684 ? 14'd14173 : 6576))) >> 3) >> 3);
            
            4'd12: result_0149 = (b * ((((a - 14'd5570) ^ (14'd1026 + a)) - ((14'd8929 ^ 14'd10105) | (b ? 14'd12812 : 2613))) ? (~b) : 12460));
            
            4'd13: result_0149 = ((b + 14'd6308) ^ 14'd11268);
            
            default: result_0149 = 14'd15932;
        endcase
    end

endmodule
        