
module simple_alu_0291(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0291
);

    always @(*) begin
        case(op)
            
            4'd0: result_0291 = ((a ^ b) ^ ((~(14'd11761 + (14'd15035 << 1))) >> 2));
            
            4'd1: result_0291 = (((14'd12248 - (14'd3888 >> 3)) << 1) + (~((14'd12835 ? (14'd3646 >> 3) : 6898) + ((a + b) | (14'd7919 - 14'd2048)))));
            
            4'd2: result_0291 = ((b + 14'd13797) - (b >> 2));
            
            4'd3: result_0291 = (14'd1683 ^ (~((14'd13365 ^ (b - 14'd8863)) & ((b ^ 14'd14595) - (14'd6561 * b)))));
            
            4'd4: result_0291 = ((~(((b ? b : 1141) << 3) * a)) ? (14'd16349 << 1) : 10324);
            
            4'd5: result_0291 = (~14'd4639);
            
            4'd6: result_0291 = (((a & b) >> 1) ^ ((14'd300 & ((14'd7945 - b) >> 2)) ^ (((14'd11335 | a) - 14'd163) ^ ((~14'd1109) ? a : 13611))));
            
            4'd7: result_0291 = (~((a - ((14'd10359 << 1) ^ (~a))) - (14'd5933 - ((14'd8818 - b) ^ (14'd5138 ? a : 8022)))));
            
            4'd8: result_0291 = (14'd12144 >> 1);
            
            4'd9: result_0291 = (~14'd5626);
            
            4'd10: result_0291 = (((~(a ^ (14'd2128 >> 3))) + (b * ((14'd11157 ^ 14'd7140) ? (14'd12427 - 14'd9284) : 8164))) ? ((((a | a) | (a ? a : 8552)) - a) | a) : 5746);
            
            4'd11: result_0291 = (~(((14'd3623 + (14'd8863 >> 2)) << 2) ^ b));
            
            4'd12: result_0291 = (((14'd11581 & (14'd3370 ? b : 14080)) | (((b & 14'd4184) ^ (b >> 1)) << 3)) + ((((b | 14'd7342) ^ (14'd12073 + b)) + 14'd13680) & (14'd9048 ^ (~(14'd8467 | 14'd9983)))));
            
            default: result_0291 = 14'd1109;
        endcase
    end

endmodule
        