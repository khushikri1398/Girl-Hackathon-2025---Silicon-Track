
module simple_alu_0070(
    input [11:0] a, b,
    input [3:0] op,
    output reg [11:0] result_0070
);

    always @(*) begin
        case(op)
            
            4'd0: result_0070 = ((((~12'd3678) ? (12'd3500 - 12'd4054) : 3862) ? ((b + b) ^ (12'd2183 - b)) : 2614) - (((12'd1750 - a) & (a ? b : 2781)) - 12'd2759));
            
            4'd1: result_0070 = ((((b << 2) + (~12'd2204)) * (a ^ (12'd166 | 12'd2336))) ^ (((~12'd3354) >> 3) * ((12'd2979 * 12'd2843) - (~12'd2301))));
            
            4'd2: result_0070 = (~(((12'd2353 << 2) - (b - a)) - ((12'd3308 >> 2) * (b ? b : 447))));
            
            4'd3: result_0070 = (a >> 1);
            
            4'd4: result_0070 = ((12'd4071 | (12'd1579 ^ (~b))) + 12'd1624);
            
            4'd5: result_0070 = ((~((12'd2076 * 12'd4012) + (a >> 2))) ^ b);
            
            4'd6: result_0070 = ((((12'd2393 - 12'd540) * 12'd2592) - ((~12'd2882) ? (a | 12'd2002) : 3262)) & ((12'd1706 | 12'd3248) ^ ((12'd933 * b) ? (b >> 3) : 3031)));
            
            4'd7: result_0070 = ((12'd2632 ^ ((12'd1199 | b) + (b << 3))) | (((b + b) >> 3) - ((~12'd108) - (a * b))));
            
            4'd8: result_0070 = ((12'd1284 & ((~12'd1633) & (12'd2567 ^ b))) & (((12'd16 + 12'd3887) ? (b ^ a) : 2087) + (12'd3589 * (a | 12'd2223))));
            
            4'd9: result_0070 = ((((a + a) | (12'd2045 - b)) ? 12'd3922 : 1527) | (((12'd1914 | 12'd3070) << 3) << 2));
            
            4'd10: result_0070 = ((12'd2815 + ((12'd1324 | 12'd906) ^ (12'd3285 | 12'd3798))) + a);
            
            4'd11: result_0070 = ((((b << 1) & (b << 3)) | a) | b);
            
            4'd12: result_0070 = (12'd3085 & 12'd2816);
            
            4'd13: result_0070 = ((12'd1896 + (12'd1311 ? (a + 12'd810) : 3400)) + (a + 12'd184));
            
            default: result_0070 = b;
        endcase
    end

endmodule
        