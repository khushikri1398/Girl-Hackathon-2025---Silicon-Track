
module simple_alu_0863(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0863
);

    always @(*) begin
        case(op)
            
            4'd0: result_0863 = (((14'd4775 >> 1) | (14'd9494 - 14'd9059)) ^ ((((14'd3698 ? 14'd12397 : 4962) << 3) + ((14'd14640 ^ b) ^ (~14'd12514))) >> 3));
            
            4'd1: result_0863 = (b ^ ((14'd5772 + ((b | a) - 14'd14935)) >> 2));
            
            4'd2: result_0863 = (((((a ^ a) ^ (a & b)) & 14'd13749) & (((a & 14'd15772) * (14'd4305 ^ 14'd3299)) & ((14'd9778 >> 3) & (b ^ 14'd13219)))) ^ ((14'd2512 ^ (~(a ^ a))) - (((a ^ 14'd8410) | (14'd682 ^ 14'd10253)) << 2)));
            
            default: result_0863 = 14'd8828;
        endcase
    end

endmodule
        