
module simple_alu_0015(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0015
);

    always @(*) begin
        case(op)
            
            4'd0: result_0015 = (((((14'd9409 ? 14'd675 : 16150) - 14'd4009) + ((14'd11782 ? a : 5705) - (~14'd11372))) << 1) ? ((((14'd10256 - b) ^ (b | b)) << 3) - (((b * a) & (a * 14'd5532)) ^ ((14'd10590 * 14'd6180) - 14'd4806))) : 6375);
            
            4'd1: result_0015 = ((b + (a & (b * 14'd2742))) & (((~(14'd13966 & 14'd15832)) ? ((14'd10173 ^ a) - (a ? 14'd16113 : 8644)) : 827) | ((14'd2487 * b) << 1)));
            
            4'd2: result_0015 = (~((~((b ? b : 5672) + (14'd8026 << 1))) << 3));
            
            4'd3: result_0015 = ((((14'd873 & 14'd14387) ^ (14'd9434 - (14'd11759 << 3))) ? ((b >> 1) << 3) : 16119) - ((~(14'd3892 * 14'd9735)) - (((b - 14'd13538) + (14'd7678 ^ 14'd13565)) | (14'd3113 | (14'd3386 + a)))));
            
            4'd4: result_0015 = (((14'd12526 >> 3) + 14'd8371) ? ((((14'd375 & a) * (a - a)) ^ ((14'd8244 ? b : 4853) ? (14'd7744 << 1) : 1129)) >> 2) : 8359);
            
            4'd5: result_0015 = (((14'd14035 ^ ((14'd8534 | 14'd4430) * (a + 14'd4098))) & a) | 14'd13177);
            
            4'd6: result_0015 = (((14'd12760 ? ((a << 1) * 14'd5634) : 11065) ^ ((14'd7588 * 14'd13905) ^ (14'd9808 & (a >> 3)))) + ((((~14'd6063) ? (b | a) : 10649) & ((14'd16364 ^ b) << 1)) | (14'd6604 << 1)));
            
            4'd7: result_0015 = ((14'd940 | (((14'd12726 ^ 14'd14319) * (~a)) | ((~a) - 14'd10973))) ? ((a | 14'd5084) >> 3) : 5832);
            
            4'd8: result_0015 = ((((14'd15694 - 14'd3635) + (~(14'd2118 << 1))) - (((14'd263 - 14'd9945) * (b ? a : 995)) + (b & (a & b)))) + (14'd13384 << 1));
            
            4'd9: result_0015 = ((14'd11427 & (~(~(b + 14'd4016)))) ? ((((b ? b : 14708) & (a << 3)) + ((~14'd12388) | (b & b))) * (14'd12265 << 2)) : 9725);
            
            4'd10: result_0015 = ((14'd4556 * (((14'd3367 >> 2) ? (a ^ 14'd5794) : 10212) ^ ((a - b) << 3))) ^ ((((14'd8750 >> 1) & 14'd7393) >> 3) + ((~(14'd4947 * b)) & ((b ? 14'd9340 : 12578) & (14'd14562 + 14'd15342)))));
            
            4'd11: result_0015 = ((((b + (14'd3879 ? a : 9003)) >> 3) >> 1) >> 1);
            
            4'd12: result_0015 = (((~((b ^ 14'd15611) | a)) + (((14'd15273 + b) ? (b - 14'd11163) : 11950) ? ((a + a) >> 2) : 13707)) - ((14'd529 * (b << 1)) ? 14'd10179 : 2309));
            
            4'd13: result_0015 = (b * (14'd1406 ? (((14'd15790 ? b : 8018) >> 1) >> 2) : 12661));
            
            4'd14: result_0015 = (((((b - 14'd1439) ^ (14'd1984 & a)) * a) ^ a) ? 14'd3908 : 7133);
            
            4'd15: result_0015 = ((b * (a & ((~b) - (14'd15979 >> 1)))) ^ ((~(b * 14'd13699)) << 1));
            
            default: result_0015 = a;
        endcase
    end

endmodule
        