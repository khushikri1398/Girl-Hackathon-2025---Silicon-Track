
module simple_alu_0071(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0071
);

    always @(*) begin
        case(op)
            
            4'd0: result_0071 = ((14'd3791 * (b + ((14'd8494 << 3) | (14'd5751 | 14'd14583)))) ^ ((a + 14'd8311) << 1));
            
            4'd1: result_0071 = (14'd6180 ^ ((((14'd12870 << 1) ^ a) & (~(~b))) * ((b ^ (a ? a : 6065)) * ((~14'd13887) & (~14'd14596)))));
            
            4'd2: result_0071 = ((~(~14'd8743)) + a);
            
            4'd3: result_0071 = ((~(~(~(14'd12402 >> 1)))) - (b << 1));
            
            4'd4: result_0071 = (~(((14'd2651 & (a - b)) - 14'd4209) & ((14'd4893 >> 3) >> 2)));
            
            4'd5: result_0071 = ((~(((14'd670 << 2) >> 3) ? ((14'd16130 ? b : 1984) >> 3) : 12348)) * ((b - ((b & b) << 3)) ? 14'd9866 : 7852));
            
            4'd6: result_0071 = ((((a << 1) - (a ? b : 13708)) - b) << 1);
            
            default: result_0071 = a;
        endcase
    end

endmodule
        