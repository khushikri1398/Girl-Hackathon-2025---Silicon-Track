
module pipeline_0520(
    input clk,
    input rst_n,
    input [5:0] data_in,
    input [1:0] control,
    output reg [5:0] result_0520
);

    // Pipeline registers
    
    reg [5:0] stage0_reg;
    wire [5:0] stage0_next;
    
    reg [5:0] stage1_reg;
    wire [5:0] stage1_next;
    
    reg [5:0] stage2_reg;
    wire [5:0] stage2_next;
    
    
    // Combinational logic for each stage
    
    
    assign stage0_next = data_in;
    
    
    
    assign stage1_next = stage0_reg;
    
    
    
    assign stage2_next = stage1_reg;
    
    
    
    // Pipeline registers update
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            
            stage0_reg <= 6'd0;
            
            stage1_reg <= 6'd0;
            
            stage2_reg <= 6'd0;
            
        end else begin
            
            
            stage0_reg <= stage0_next;
            
            
            
            stage1_reg <= stage1_next;
            
            
            
            stage2_reg <= stage2_next;
            
            
        end
    end
    
    // Output selection based on control
    always @(*) begin
        case(control)
            
            2'd0: result_0520 = stage0_reg;
            
            2'd1: result_0520 = stage1_reg;
            
            2'd2: result_0520 = stage2_reg;
            
            default: result_0520 = stage2_reg;
        endcase
    end

endmodule
        