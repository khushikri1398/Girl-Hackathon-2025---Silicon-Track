
module simple_alu_0972(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0972
);

    always @(*) begin
        case(op)
            
            4'd0: result_0972 = (((((14'd13976 + 14'd11941) ^ (14'd2464 - a)) >> 2) ? (((14'd4081 ? b : 5801) ^ (a ? 14'd399 : 3722)) + b) : 11212) | 14'd5207);
            
            4'd1: result_0972 = (14'd12324 * (14'd1992 + 14'd2347));
            
            4'd2: result_0972 = ((~14'd15948) << 3);
            
            4'd3: result_0972 = ((14'd12887 + ((~(b ? 14'd14134 : 13985)) ^ (~(a ^ 14'd11402)))) << 2);
            
            4'd4: result_0972 = (((((14'd7723 ^ 14'd11233) * (14'd13656 << 2)) ^ ((14'd2138 ^ 14'd15959) ? (~14'd11970) : 15580)) * (14'd427 - ((14'd10766 * 14'd7083) & (14'd391 * 14'd10138)))) >> 3);
            
            4'd5: result_0972 = (14'd11087 + (((~(14'd9874 >> 2)) | ((14'd9106 & 14'd2712) >> 3)) - 14'd4799));
            
            4'd6: result_0972 = (((14'd8141 >> 1) << 2) ^ b);
            
            4'd7: result_0972 = (14'd2283 * a);
            
            4'd8: result_0972 = (a & 14'd6808);
            
            4'd9: result_0972 = (14'd14362 << 3);
            
            4'd10: result_0972 = (a & ((14'd10877 ^ 14'd13261) * 14'd6857));
            
            4'd11: result_0972 = ((14'd249 & (((14'd4423 << 2) * (b * 14'd15117)) * 14'd3460)) ^ (b >> 2));
            
            4'd12: result_0972 = (~14'd15451);
            
            4'd13: result_0972 = (((b & ((~a) >> 1)) & (14'd15361 * 14'd8876)) << 1);
            
            default: result_0972 = 14'd2000;
        endcase
    end

endmodule
        