
module simple_alu_0074(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0074
);

    always @(*) begin
        case(op)
            
            4'd0: result_0074 = (a ? (~b) : 9781);
            
            4'd1: result_0074 = (((14'd6454 >> 2) & (((b ^ 14'd14241) * 14'd13376) & (a << 1))) >> 3);
            
            4'd2: result_0074 = ((a ? ((14'd3470 ^ (14'd5708 + b)) << 3) : 9280) << 2);
            
            4'd3: result_0074 = (14'd6177 ^ 14'd7583);
            
            4'd4: result_0074 = (~(((~(14'd10432 ^ 14'd7127)) | ((~b) ? (14'd194 - 14'd2403) : 6427)) >> 2));
            
            4'd5: result_0074 = (~((b << 1) & (((14'd1778 - b) | (14'd15992 << 3)) - ((b & 14'd9956) | (14'd16233 * 14'd15427)))));
            
            4'd6: result_0074 = (a - (((14'd9879 * (~14'd7354)) | ((14'd9514 ^ 14'd13325) >> 1)) * ((a & (14'd2858 + a)) - b)));
            
            4'd7: result_0074 = (a | ((((a >> 2) >> 1) ? a : 1937) >> 3));
            
            4'd8: result_0074 = (((((~14'd12770) & (~14'd9335)) | ((b << 1) << 1)) >> 3) & (~(b * (14'd1336 | (14'd13655 ^ 14'd1404)))));
            
            4'd9: result_0074 = (14'd11306 ^ ((((a >> 1) ? (b | 14'd2715) : 8555) ^ (~(14'd3362 + 14'd15887))) | (14'd5252 << 2)));
            
            4'd10: result_0074 = ((((14'd8958 - (14'd15478 & a)) << 1) & 14'd45) >> 2);
            
            default: result_0074 = b;
        endcase
    end

endmodule
        