
module simple_alu_0921(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0921
);

    always @(*) begin
        case(op)
            
            4'd0: result_0921 = (((((14'd13975 + a) ^ (14'd12906 >> 1)) - a) ? (((14'd14348 - 14'd10949) & b) ? (14'd8965 << 1) : 13735) : 7032) << 1);
            
            4'd1: result_0921 = ((((~14'd13279) + ((b * 14'd3834) & (a >> 2))) | (((b ? 14'd9433 : 8523) | (b & 14'd6137)) << 3)) * ((14'd2703 ? ((14'd744 ? a : 10293) * 14'd15021) : 15084) << 1));
            
            4'd2: result_0921 = (b ? ((((14'd14005 ? 14'd8551 : 9121) ^ (~14'd9885)) | ((14'd11222 << 2) + (~14'd13508))) >> 1) : 10158);
            
            4'd3: result_0921 = (14'd4957 + (((~(b >> 3)) >> 2) * b));
            
            4'd4: result_0921 = (((b ? (14'd15640 | (b + b)) : 4228) ? b : 4290) * ((b << 2) ? 14'd237 : 10440));
            
            4'd5: result_0921 = ((14'd8334 & a) ? (a ^ (((a ? 14'd13747 : 14444) & (14'd11621 >> 3)) + (~a))) : 6691);
            
            4'd6: result_0921 = (((((14'd5226 | 14'd10185) + (14'd8727 - 14'd14242)) * 14'd8720) + a) << 2);
            
            4'd7: result_0921 = (((14'd1015 & ((a << 3) ^ (14'd10760 ^ 14'd1836))) ^ 14'd7425) & ((((14'd7153 - 14'd6941) - (b + a)) - (~(14'd4513 | 14'd551))) | (((a << 2) ^ (14'd9363 | a)) ^ b)));
            
            4'd8: result_0921 = ((14'd15391 & (((14'd3753 ^ b) << 2) + (14'd5057 & (a | b)))) | 14'd9079);
            
            4'd9: result_0921 = (~(a << 1));
            
            4'd10: result_0921 = (a | ((14'd14290 - ((~14'd13075) * 14'd16101)) | ((14'd12651 | 14'd6276) & ((14'd1325 * 14'd8427) >> 3))));
            
            4'd11: result_0921 = (((14'd5920 + ((14'd11566 + 14'd12469) + 14'd13606)) | (14'd13431 * (~(a << 2)))) + 14'd15522);
            
            4'd12: result_0921 = (((((~14'd8077) >> 2) >> 2) ^ (((14'd2029 + 14'd43) << 1) | 14'd2778)) ^ b);
            
            default: result_0921 = a;
        endcase
    end

endmodule
        