
module simple_alu_0108(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0108
);

    always @(*) begin
        case(op)
            
            4'd0: result_0108 = (((((b ? 14'd9040 : 70) | (a >> 2)) ? b : 7385) ? ((~(14'd3908 << 3)) >> 3) : 2540) ? (14'd3639 ? (((14'd6669 >> 2) * 14'd14845) + ((14'd2529 - a) ? 14'd13397 : 13479)) : 10097) : 15536);
            
            4'd1: result_0108 = ((14'd5256 + (((14'd13434 | 14'd6892) >> 2) * 14'd7772)) << 2);
            
            4'd2: result_0108 = (14'd16087 << 3);
            
            4'd3: result_0108 = ((14'd8162 - (((14'd3988 + a) - (a >> 1)) << 3)) ? (((~(a | 14'd10090)) - ((~14'd15602) ^ (14'd13636 ? 14'd3858 : 2462))) + ((a ^ (b ^ 14'd485)) | (~14'd10190))) : 8321);
            
            4'd4: result_0108 = (((((a << 3) * (14'd1398 >> 1)) & ((a | 14'd10558) + (14'd6592 * 14'd13276))) >> 1) | ((14'd11574 | (14'd480 * (b >> 3))) | (((a + a) & (14'd10381 ^ b)) ^ ((14'd13123 - a) << 2))));
            
            4'd5: result_0108 = (((a | a) | (((14'd15748 - a) ^ (14'd13755 << 3)) & a)) ? b : 16186);
            
            4'd6: result_0108 = ((~(14'd859 - (b << 2))) >> 3);
            
            4'd7: result_0108 = ((((14'd12646 * (~14'd3746)) >> 1) + (((a ^ b) + (a & 14'd16063)) >> 3)) >> 1);
            
            4'd8: result_0108 = ((14'd10920 << 3) >> 3);
            
            4'd9: result_0108 = ((~14'd12489) ? ((b | ((14'd7225 + 14'd1621) | (14'd14124 * 14'd10068))) ? (((a & 14'd5366) >> 2) - ((b * b) >> 2)) : 6536) : 14214);
            
            4'd10: result_0108 = (((((b - 14'd12659) - 14'd14477) * ((a ? a : 7835) | (14'd7754 & 14'd8497))) ^ 14'd8152) + 14'd10711);
            
            4'd11: result_0108 = ((b + b) >> 1);
            
            4'd12: result_0108 = (((b + 14'd9330) + (~((a * a) | (a - b)))) >> 1);
            
            default: result_0108 = a;
        endcase
    end

endmodule
        