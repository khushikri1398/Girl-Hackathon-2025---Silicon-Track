
module simple_alu_0322(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0322
);

    always @(*) begin
        case(op)
            
            4'd0: result_0322 = (((((14'd256 + 14'd10613) & 14'd7560) | (~(b ^ b))) + (a + 14'd9952)) << 1);
            
            4'd1: result_0322 = (((((14'd7919 & 14'd14672) ? 14'd15843 : 6849) | ((~14'd6772) & (14'd1818 - a))) >> 2) | (a | ((14'd1489 + a) & (~(14'd201 - 14'd2806)))));
            
            4'd2: result_0322 = (((~(a ^ (14'd15883 << 1))) | (14'd10878 * ((14'd9800 + 14'd567) << 1))) + ((14'd7272 | 14'd5199) >> 2));
            
            4'd3: result_0322 = (((((14'd3376 & 14'd1351) * (a * 14'd7511)) + ((14'd4029 ? 14'd15969 : 11723) ? (14'd245 + a) : 15122)) & (((~14'd13053) << 2) ^ (14'd9061 - 14'd6669))) ^ (((14'd15715 - 14'd1297) & 14'd13418) >> 3));
            
            4'd4: result_0322 = (14'd1741 - b);
            
            4'd5: result_0322 = ((~b) - (((~b) ? ((14'd12429 << 2) >> 1) : 6034) & (((14'd9729 ^ 14'd16043) >> 1) & (14'd14765 * (14'd5652 - b)))));
            
            4'd6: result_0322 = (14'd15081 << 1);
            
            4'd7: result_0322 = (b & (~(((14'd4075 + b) << 2) ? (b * 14'd4855) : 14700)));
            
            4'd8: result_0322 = (14'd12007 ^ (((~b) ? ((14'd4879 & b) << 3) : 15118) + (((14'd14413 ? 14'd8991 : 1399) - (14'd9267 * 14'd3008)) | ((14'd5803 ? 14'd5519 : 14883) & (14'd14088 & b)))));
            
            4'd9: result_0322 = ((b | ((14'd11682 << 1) + ((14'd3055 >> 2) ? (14'd2001 >> 1) : 2518))) ? 14'd1988 : 9404);
            
            4'd10: result_0322 = ((~14'd8429) ^ ((b | 14'd15029) & ((14'd1194 << 3) ? (~(b & 14'd4654)) : 15233)));
            
            4'd11: result_0322 = (((14'd8895 ? ((14'd12495 ? a : 10255) | 14'd10825) : 8317) * (((14'd6026 ^ 14'd3389) * b) ^ ((b & a) * a))) << 1);
            
            4'd12: result_0322 = (((~((14'd4215 - 14'd11728) >> 1)) ^ (((14'd558 + 14'd5601) ^ b) ? 14'd2765 : 12894)) & (((~(a & 14'd14812)) ^ 14'd11782) << 1));
            
            4'd13: result_0322 = (~14'd8061);
            
            4'd14: result_0322 = (((((a + 14'd14693) ^ (~14'd7006)) - ((a << 2) ^ (14'd1357 + a))) & (((b - a) | (a ? 14'd7456 : 6769)) | 14'd9752)) | ((((14'd13048 >> 1) >> 3) >> 3) & ((~(14'd5 - 14'd9490)) ? ((14'd15915 & a) ? a : 12961) : 7634)));
            
            default: result_0322 = a;
        endcase
    end

endmodule
        