
module simple_alu_0748(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0748
);

    always @(*) begin
        case(op)
            
            4'd0: result_0748 = ((((~(14'd9273 * 14'd3865)) & ((14'd3488 ? 14'd10970 : 2225) << 2)) ^ (14'd7540 | (b * (~a)))) * ((14'd10238 * ((14'd9724 + b) ^ (14'd12588 & 14'd28))) | (14'd5908 | ((a & 14'd2479) >> 3))));
            
            4'd1: result_0748 = ((14'd2758 - (((14'd16205 >> 1) & b) << 1)) | a);
            
            4'd2: result_0748 = ((((14'd5565 * (a << 1)) | ((14'd14379 & a) >> 2)) ? ((14'd7990 ^ (~14'd93)) | ((14'd13698 ^ 14'd10726) >> 1)) : 15733) | ((~((14'd3136 + 14'd13402) | (14'd8479 | a))) << 3));
            
            4'd3: result_0748 = (14'd3340 | b);
            
            4'd4: result_0748 = (14'd146 >> 2);
            
            4'd5: result_0748 = (((14'd10000 - 14'd7675) - b) & ((((14'd14934 >> 2) ? (a ? 14'd15715 : 4859) : 8021) & ((14'd12648 - 14'd15814) & (14'd4453 ^ 14'd1780))) ^ (((b & 14'd15052) + 14'd96) ^ 14'd7720)));
            
            4'd6: result_0748 = (((a ^ 14'd900) | ((~14'd10862) << 3)) ^ a);
            
            4'd7: result_0748 = ((((14'd539 * (b << 3)) << 2) >> 3) + (14'd12948 * (((b | 14'd10804) - (a >> 2)) << 2)));
            
            default: result_0748 = 14'd10062;
        endcase
    end

endmodule
        