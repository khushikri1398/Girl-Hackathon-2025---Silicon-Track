
module simple_alu_0089(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0089
);

    always @(*) begin
        case(op)
            
            4'd0: result_0089 = (((((14'd15972 * a) << 3) + 14'd15903) & (~((a ? 14'd8581 : 9146) ? (14'd14396 - a) : 15214))) << 2);
            
            4'd1: result_0089 = (~((b << 2) >> 1));
            
            4'd2: result_0089 = (a * ((((14'd15600 ^ a) & 14'd15159) + ((14'd12456 + a) | (14'd1294 >> 1))) ^ (((b | b) & b) << 2)));
            
            4'd3: result_0089 = ((((b << 1) >> 3) >> 3) ? (((~14'd5031) ? ((a & 14'd11899) >> 2) : 6565) << 2) : 16013);
            
            4'd4: result_0089 = ((a ^ (14'd1286 | (a << 3))) + (a * (b & a)));
            
            4'd5: result_0089 = ((~(~((a * 14'd11444) << 2))) ^ ((((14'd13750 ^ a) ^ (a * b)) ? (14'd5260 + (14'd13843 & b)) : 11487) - (~(~(a | 14'd16217)))));
            
            4'd6: result_0089 = ((a * b) | ((((14'd1187 + 14'd3411) >> 1) * 14'd11321) >> 2));
            
            4'd7: result_0089 = (((14'd7966 | ((14'd892 ? b : 11628) ^ (a ^ a))) & (((a ^ b) * (b & 14'd16243)) ? ((b & 14'd14928) * a) : 8390)) ^ ((((14'd8767 - a) ? (14'd8482 & b) : 11550) >> 3) + (a << 2)));
            
            4'd8: result_0089 = ((14'd15437 - 14'd12689) ^ (~a));
            
            4'd9: result_0089 = ((((~b) & ((14'd8779 + a) << 1)) ? 14'd3812 : 584) - (14'd6536 ? (((b ^ a) ? (~b) : 13135) << 2) : 13128));
            
            4'd10: result_0089 = ((((14'd11759 << 1) & ((~b) ^ (14'd7389 + 14'd9218))) | (((14'd3561 * 14'd10726) + 14'd9843) << 2)) >> 2);
            
            4'd11: result_0089 = (14'd15506 - ((((14'd14267 & b) & (a << 3)) >> 1) << 1));
            
            4'd12: result_0089 = ((14'd15470 ? (((14'd6931 - 14'd6392) - 14'd12773) + ((b ? 14'd5844 : 2285) ^ (14'd1381 + 14'd10769))) : 13111) ^ (((~(a << 2)) & a) - (~14'd14823)));
            
            4'd13: result_0089 = (b ^ (~(a >> 3)));
            
            4'd14: result_0089 = (14'd11549 | (14'd2894 & (b * ((~b) << 1))));
            
            default: result_0089 = a;
        endcase
    end

endmodule
        