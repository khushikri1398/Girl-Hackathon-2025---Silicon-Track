
module simple_alu_0013(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0013
);

    always @(*) begin
        case(op)
            
            4'd0: result_0013 = (b >> 1);
            
            4'd1: result_0013 = (((~((14'd4263 ? b : 7958) ? 14'd11200 : 7094)) + (((14'd187 & 14'd14152) & (14'd368 + a)) | ((a & 14'd6339) + (b << 2)))) ? (~(((b >> 2) | (14'd546 ^ b)) * ((14'd5043 >> 1) & (14'd3094 + a)))) : 9462);
            
            4'd2: result_0013 = ((a << 3) >> 2);
            
            4'd3: result_0013 = (((((14'd3633 & 14'd15394) + b) ^ ((~14'd6102) >> 1)) * (((a & a) + (14'd12876 + 14'd11375)) - ((14'd1426 << 3) ? (a >> 1) : 3321))) << 1);
            
            4'd4: result_0013 = (((~((b ? 14'd5628 : 13426) + (~14'd12386))) * (b << 2)) * ((14'd1574 + (~(a + 14'd7062))) - ((b * (b - 14'd4926)) << 2)));
            
            4'd5: result_0013 = (((((14'd11021 * 14'd10566) << 2) ^ ((14'd3633 | b) * 14'd11280)) * (((b + 14'd5055) ? (~14'd9134) : 4058) & (a << 1))) >> 2);
            
            4'd6: result_0013 = (((~((a >> 1) ^ (14'd12863 ^ 14'd5490))) & (((a << 1) ^ (14'd11440 << 3)) << 3)) << 1);
            
            4'd7: result_0013 = (~(14'd2998 * 14'd235));
            
            4'd8: result_0013 = (14'd3330 ^ ((14'd15633 * ((14'd12435 ^ a) >> 1)) - ((14'd15728 >> 1) | 14'd883)));
            
            4'd9: result_0013 = ((14'd11854 - (b - 14'd646)) + ((((a >> 1) | (b ? 14'd13634 : 7858)) << 2) - (((a >> 3) ^ (b ? 14'd5802 : 874)) << 3)));
            
            4'd10: result_0013 = ((a + (((14'd10503 ? a : 11540) & (14'd14439 ^ 14'd9538)) - (~14'd628))) << 1);
            
            4'd11: result_0013 = ((((~(14'd8919 * b)) * (14'd37 ^ (14'd14840 ? 14'd16326 : 14126))) & (14'd14034 & ((a * b) >> 2))) ? (14'd11770 >> 1) : 3651);
            
            default: result_0013 = b;
        endcase
    end

endmodule
        