
module simple_alu_0876(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0876
);

    always @(*) begin
        case(op)
            
            4'd0: result_0876 = (((((b ^ 14'd10002) ^ (14'd8991 - 14'd8915)) & (~(b - 14'd14247))) ^ (((b - 14'd15114) - (b << 3)) ? (b - (a * 14'd748)) : 2151)) + 14'd300);
            
            4'd1: result_0876 = (b - 14'd183);
            
            4'd2: result_0876 = ((((14'd10030 & 14'd1371) >> 1) + (a ^ 14'd7254)) | (b & 14'd6074));
            
            4'd3: result_0876 = (((((14'd3215 - a) ^ a) + 14'd14617) - 14'd14210) | ((((14'd6709 ? b : 5018) ? (14'd4357 ? a : 7904) : 15980) >> 2) >> 2));
            
            4'd4: result_0876 = (~14'd12781);
            
            4'd5: result_0876 = (((((a | 14'd11158) & (14'd598 ? 14'd14219 : 12978)) >> 3) | (((a << 2) - 14'd3389) ^ ((14'd12394 << 3) - (~a)))) >> 2);
            
            4'd6: result_0876 = (14'd15225 + a);
            
            4'd7: result_0876 = (14'd5621 ^ a);
            
            4'd8: result_0876 = (((~((14'd12965 | 14'd7467) << 1)) >> 1) - (b - (~((14'd9856 >> 1) ? (a + b) : 1627))));
            
            4'd9: result_0876 = ((((~(a & 14'd3403)) * (14'd1507 + (~14'd69))) * b) & (~a));
            
            4'd10: result_0876 = (14'd13437 - (a + (((b + 14'd11975) + a) ^ (14'd8449 - (b >> 3)))));
            
            4'd11: result_0876 = (((((b * a) + (14'd15436 >> 3)) >> 2) + (((14'd15617 << 1) - (14'd12604 ? a : 2606)) - 14'd4899)) * (14'd9679 >> 2));
            
            4'd12: result_0876 = (((b >> 1) * 14'd2385) << 3);
            
            4'd13: result_0876 = ((14'd4621 & ((14'd3273 * b) | (14'd15352 ^ (14'd9889 & a)))) << 3);
            
            4'd14: result_0876 = ((a >> 3) & a);
            
            default: result_0876 = a;
        endcase
    end

endmodule
        