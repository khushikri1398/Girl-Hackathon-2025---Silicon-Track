
module simple_alu_0145(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0145
);

    always @(*) begin
        case(op)
            
            4'd0: result_0145 = (14'd5562 << 2);
            
            4'd1: result_0145 = ((((a >> 2) + (14'd531 - (~14'd3870))) + 14'd9728) + (14'd2898 ? (14'd11822 + (14'd3544 | (14'd925 & 14'd9107))) : 9430));
            
            4'd2: result_0145 = ((((14'd10399 * (a << 1)) & ((14'd9567 ? 14'd10789 : 4470) << 2)) | (((14'd4827 ? 14'd9057 : 10480) ^ 14'd5924) * ((a & 14'd2660) ^ (a * 14'd9545)))) & (a + 14'd7174));
            
            4'd3: result_0145 = (((((14'd8153 ^ b) ? (14'd11563 * 14'd5007) : 12039) ? (b ? (b ^ b) : 10670) : 13734) + (a << 2)) | (14'd4760 | ((~(14'd12416 ? 14'd16328 : 9408)) * a)));
            
            4'd4: result_0145 = (a ? (a * ((14'd6716 - a) * 14'd205)) : 13682);
            
            4'd5: result_0145 = (b ? (((~(14'd4068 * a)) << 1) << 1) : 3152);
            
            4'd6: result_0145 = (((14'd11281 ? (14'd0 - (14'd6400 & 14'd13170)) : 15739) - (14'd2085 + (14'd7463 >> 1))) & 14'd13493);
            
            4'd7: result_0145 = (14'd2126 & (~(14'd14626 >> 1)));
            
            4'd8: result_0145 = (((~((b - 14'd14828) & (14'd3500 + b))) << 2) - (14'd14179 << 3));
            
            default: result_0145 = 14'd14568;
        endcase
    end

endmodule
        