
module simple_alu_0258(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0258
);

    always @(*) begin
        case(op)
            
            4'd0: result_0258 = ((a - (((14'd9699 - 14'd13585) << 1) << 3)) | 14'd3773);
            
            4'd1: result_0258 = ((((a >> 3) - 14'd3380) * 14'd6363) & 14'd4076);
            
            4'd2: result_0258 = ((14'd11065 + 14'd10076) - (((14'd10052 ? 14'd10671 : 11274) ^ b) & 14'd575));
            
            4'd3: result_0258 = (((((14'd12466 - a) - (14'd16051 - 14'd4746)) >> 3) * (b ^ ((a >> 3) * 14'd14340))) ? b : 16220);
            
            4'd4: result_0258 = (((~a) << 2) * ((((b >> 2) + b) ? ((~a) | 14'd9783) : 5529) + b));
            
            4'd5: result_0258 = ((14'd10189 ^ (((14'd8880 ? 14'd11240 : 3137) >> 2) ^ (~(a ? b : 1353)))) << 3);
            
            4'd6: result_0258 = (14'd7851 << 1);
            
            4'd7: result_0258 = (((14'd10507 | (b ? 14'd5554 : 8200)) + 14'd2712) ? (~(14'd12920 * a)) : 2862);
            
            4'd8: result_0258 = ((a << 1) ^ 14'd3738);
            
            4'd9: result_0258 = (~((~b) - ((14'd11731 | a) * ((b & 14'd16363) << 3))));
            
            4'd10: result_0258 = ((((14'd16163 + (~b)) - ((14'd4874 ^ b) >> 1)) << 1) >> 3);
            
            4'd11: result_0258 = (14'd9866 + ((~((14'd4056 - 14'd12187) - (14'd16232 ^ b))) & (((~a) + 14'd6387) ^ ((14'd6485 * a) | (14'd801 >> 2)))));
            
            4'd12: result_0258 = (a ^ 14'd6459);
            
            default: result_0258 = 14'd6587;
        endcase
    end

endmodule
        