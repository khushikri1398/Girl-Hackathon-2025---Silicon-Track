
module simple_alu_0079(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0079
);

    always @(*) begin
        case(op)
            
            4'd0: result_0079 = ((~(b | a)) - a);
            
            4'd1: result_0079 = (((((14'd7160 >> 1) ? 14'd4085 : 5408) << 1) & (a ^ ((~b) >> 2))) + (b | 14'd14929));
            
            4'd2: result_0079 = ((((14'd14660 + (14'd11699 >> 1)) * (14'd15145 - (a & 14'd12094))) - (~((14'd8260 | 14'd13828) << 1))) >> 3);
            
            4'd3: result_0079 = ((14'd10366 & ((~(14'd11470 << 3)) ? ((14'd6839 - a) ^ (~14'd2846)) : 5190)) >> 3);
            
            4'd4: result_0079 = (~(14'd11010 * a));
            
            4'd5: result_0079 = ((14'd907 * 14'd434) + (((b >> 3) ? b : 4941) * ((~(14'd10044 >> 1)) * ((b ? b : 7958) ^ b))));
            
            4'd6: result_0079 = ((b ? (((b >> 2) & 14'd2666) ? ((14'd6615 << 2) << 1) : 12441) : 4992) | a);
            
            4'd7: result_0079 = (b + 14'd10287);
            
            4'd8: result_0079 = (14'd4326 & ((b & b) * (a & (~(14'd5343 ? b : 12508)))));
            
            4'd9: result_0079 = ((b ? (b * 14'd10250) : 7841) << 2);
            
            4'd10: result_0079 = ((b | (~(14'd13581 >> 3))) * a);
            
            4'd11: result_0079 = ((~14'd945) - (14'd15579 | 14'd8945));
            
            default: result_0079 = 14'd5699;
        endcase
    end

endmodule
        