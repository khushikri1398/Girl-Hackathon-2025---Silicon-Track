
module simple_alu_0478(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0478
);

    always @(*) begin
        case(op)
            
            4'd0: result_0478 = ((14'd3278 - (((14'd15863 << 3) - 14'd8058) >> 3)) >> 1);
            
            4'd1: result_0478 = ((((14'd8676 - (14'd13685 + a)) ? b : 270) - a) << 3);
            
            4'd2: result_0478 = ((((14'd4900 ^ b) * (14'd6247 | 14'd12649)) ? (14'd4252 + (14'd11320 + (b - b))) : 4596) ^ ((14'd3450 * ((14'd7680 ? 14'd13147 : 9031) * (b * 14'd10357))) << 3));
            
            4'd3: result_0478 = (((14'd1302 & (a << 1)) << 3) & ((((b & b) + b) + ((14'd4651 << 2) & 14'd4650)) ^ (((14'd14251 - 14'd8745) ^ (14'd14974 ? 14'd656 : 10566)) >> 2)));
            
            4'd4: result_0478 = (b ^ (14'd2409 ^ (14'd3337 * ((14'd319 & b) - (b ? 14'd2234 : 7333)))));
            
            4'd5: result_0478 = (((((b + 14'd992) & (14'd14363 & 14'd6580)) ^ a) ^ (((b << 1) ^ a) * b)) >> 1);
            
            4'd6: result_0478 = ((((b * a) * ((14'd7982 | a) << 3)) | 14'd15150) >> 3);
            
            default: result_0478 = 14'd2231;
        endcase
    end

endmodule
        