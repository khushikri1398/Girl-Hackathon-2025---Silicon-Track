
module simple_alu_0362(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0362
);

    always @(*) begin
        case(op)
            
            4'd0: result_0362 = (((((b >> 1) + (14'd7867 - b)) - 14'd13931) - 14'd7462) + a);
            
            4'd1: result_0362 = ((14'd10666 - 14'd15174) | ((((~b) & (14'd48 & 14'd12888)) >> 1) | b));
            
            4'd2: result_0362 = ((((a & (14'd12181 ^ b)) ? (14'd15855 + (a | b)) : 8851) ^ (14'd2311 - ((b << 3) >> 1))) ^ (b + a));
            
            4'd3: result_0362 = (((b << 3) << 2) + ((((14'd406 & 14'd11982) ^ (14'd16324 + 14'd8506)) * ((a >> 2) * (14'd12670 - a))) | (((14'd3232 & a) | (~14'd13686)) >> 3)));
            
            4'd4: result_0362 = ((((14'd5519 ? (b & 14'd12442) : 5969) << 1) & ((~(14'd15101 >> 1)) & ((14'd788 * 14'd9253) ^ (b - 14'd12178)))) - (~(14'd9341 * (~(14'd11626 << 2)))));
            
            4'd5: result_0362 = ((14'd13335 >> 1) - (((~(a | 14'd9666)) ^ ((~14'd16326) ? 14'd8400 : 11474)) << 1));
            
            4'd6: result_0362 = (14'd7146 ^ ((((14'd5265 ? 14'd13196 : 4426) ^ b) + 14'd8163) - 14'd5451));
            
            4'd7: result_0362 = (14'd3043 + (b & (14'd1587 * ((14'd7168 >> 1) - (b | 14'd11469)))));
            
            4'd8: result_0362 = (((((a & 14'd4782) | (14'd9808 & b)) & ((b | b) - (14'd16031 ? a : 9928))) | (((~14'd12084) + b) - ((14'd3794 - b) ^ (b ^ 14'd1493)))) ^ (((14'd7429 * (~a)) | ((a - 14'd8915) + (~14'd15815))) & (((b << 1) | (b | 14'd15551)) << 1)));
            
            4'd9: result_0362 = ((((~(~b)) >> 3) ? (~14'd11283) : 6981) & a);
            
            4'd10: result_0362 = (14'd1314 - ((((b ? 14'd9846 : 2030) ? 14'd16380 : 2796) & (a | (a & b))) | (((~b) | 14'd9785) >> 3)));
            
            4'd11: result_0362 = ((14'd10710 ? ((b + (14'd501 + b)) * ((14'd2889 * a) ^ b)) : 4447) | (14'd13713 ? ((b ^ b) ? 14'd5548 : 2867) : 3484));
            
            4'd12: result_0362 = ((b ^ b) << 1);
            
            default: result_0362 = 14'd11725;
        endcase
    end

endmodule
        