
module simple_alu_0338(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0338
);

    always @(*) begin
        case(op)
            
            4'd0: result_0338 = (14'd15094 << 2);
            
            4'd1: result_0338 = ((a | (((14'd4908 - 14'd10494) >> 1) + ((a | 14'd2068) * (~b)))) >> 3);
            
            4'd2: result_0338 = ((14'd12350 | (((14'd12270 & b) >> 1) & ((a * 14'd1655) | (14'd10881 >> 3)))) + 14'd2274);
            
            4'd3: result_0338 = ((((14'd14425 ^ (a - 14'd1834)) - ((14'd14358 * a) | (14'd6276 >> 2))) * (b - (14'd11498 - b))) * ((((b | 14'd3267) * (14'd5132 * 14'd7132)) ? ((a | 14'd1034) ^ (b - b)) : 4368) ? 14'd11985 : 5033));
            
            4'd4: result_0338 = (~((14'd12000 - (~(a | b))) & 14'd13837));
            
            default: result_0338 = 14'd15541;
        endcase
    end

endmodule
        