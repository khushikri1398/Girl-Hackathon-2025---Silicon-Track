
module simple_alu_0393(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0393
);

    always @(*) begin
        case(op)
            
            4'd0: result_0393 = (14'd7589 - ((~((a + 14'd9187) & (14'd3328 ? 14'd3800 : 13868))) * a));
            
            4'd1: result_0393 = (((((b ? 14'd4059 : 773) & b) & (14'd10257 << 3)) | a) - (((a ? (a + 14'd6244) : 14216) | ((a * 14'd13174) * b)) | 14'd14051));
            
            4'd2: result_0393 = (((~(14'd6594 - (~b))) & (((14'd11766 & b) >> 3) << 3)) + b);
            
            4'd3: result_0393 = (14'd6646 ? ((((a - b) << 2) | a) - ((14'd7379 | a) | (14'd560 - (a + a)))) : 9659);
            
            4'd4: result_0393 = (((((14'd4824 | 14'd13317) ^ (14'd12041 ^ 14'd7079)) & 14'd5825) * ((a - a) | b)) ^ 14'd5318);
            
            4'd5: result_0393 = (((a - b) - (a + 14'd13780)) * 14'd429);
            
            4'd6: result_0393 = (((((14'd15247 - 14'd2658) | (a - 14'd8395)) ^ ((14'd9113 | 14'd11302) ^ 14'd4552)) | (14'd9169 >> 3)) ? (((14'd6428 >> 3) << 3) >> 2) : 12682);
            
            4'd7: result_0393 = (14'd7011 ? b : 9025);
            
            4'd8: result_0393 = ((((14'd9538 << 3) * (14'd231 ^ (a ? 14'd6228 : 115))) + (((b ^ a) | (14'd2508 | 14'd4458)) + (~(14'd9563 - 14'd6760)))) ^ ((((a * a) ^ (a - 14'd9888)) & 14'd9738) - 14'd9531));
            
            default: result_0393 = 14'd885;
        endcase
    end

endmodule
        