
module simple_alu_0878(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0878
);

    always @(*) begin
        case(op)
            
            4'd0: result_0878 = ((~(((a ^ 14'd1382) ? a : 15573) >> 1)) - ((a * ((b - 14'd2260) ? (14'd9583 | 14'd1368) : 6415)) << 2));
            
            4'd1: result_0878 = ((((a ^ 14'd12123) | (b * (14'd7989 >> 2))) | (~14'd13161)) * ((((14'd2560 ^ 14'd14737) ? (~14'd5889) : 1483) << 1) << 1));
            
            4'd2: result_0878 = ((14'd4754 & (((b ? 14'd2849 : 4477) + (~14'd4879)) + ((b & 14'd13261) * 14'd6722))) << 1);
            
            4'd3: result_0878 = ((14'd4305 ? 14'd6671 : 4709) >> 2);
            
            4'd4: result_0878 = (((~a) | ((~(~14'd7283)) - ((14'd3053 ? 14'd1691 : 12320) ? (14'd1608 | 14'd8158) : 13944))) - (14'd4968 + 14'd15971));
            
            4'd5: result_0878 = (14'd13075 >> 2);
            
            4'd6: result_0878 = (b - ((14'd11796 * ((14'd13448 & 14'd5297) >> 3)) * (((b ? 14'd8525 : 13701) ? (14'd13265 | 14'd4812) : 11283) - ((b & b) + (14'd7399 | b)))));
            
            4'd7: result_0878 = (~(b ^ 14'd14322));
            
            4'd8: result_0878 = (a ? ((a ? (14'd5289 ? (14'd14732 - 14'd4652) : 12740) : 15137) * (((a | b) >> 3) & (14'd4447 + 14'd4214))) : 8322);
            
            4'd9: result_0878 = (14'd1122 + (((b | (a << 2)) & 14'd13040) + a));
            
            4'd10: result_0878 = (14'd3651 + 14'd8410);
            
            4'd11: result_0878 = (((((b - b) >> 2) << 3) >> 3) ? 14'd9232 : 6571);
            
            default: result_0878 = b;
        endcase
    end

endmodule
        