
module simple_alu_0117(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0117
);

    always @(*) begin
        case(op)
            
            4'd0: result_0117 = (b | (14'd133 << 2));
            
            4'd1: result_0117 = (14'd3033 ? (((~(14'd2343 | a)) & 14'd16336) | (((14'd16364 >> 1) * (14'd14934 ^ 14'd4058)) >> 3)) : 4050);
            
            4'd2: result_0117 = (((~((14'd13591 & 14'd15609) | (a * 14'd15354))) ^ (((a >> 2) | (14'd9409 ^ a)) >> 1)) ^ a);
            
            4'd3: result_0117 = ((~b) + (b >> 3));
            
            4'd4: result_0117 = ((~14'd5399) ^ (b ^ (b >> 1)));
            
            4'd5: result_0117 = (a & ((~(14'd11624 ^ b)) * 14'd5963));
            
            4'd6: result_0117 = (((14'd6201 << 2) << 3) ^ 14'd11718);
            
            4'd7: result_0117 = ((14'd4774 ? ((~(b * a)) << 2) : 11977) | (~14'd6552));
            
            4'd8: result_0117 = (((((14'd8988 + 14'd5724) ^ (14'd125 >> 3)) & 14'd8463) >> 2) & (~((~(14'd7208 ? a : 15973)) - ((14'd8603 ? 14'd436 : 12180) * (14'd2857 & 14'd15353)))));
            
            4'd9: result_0117 = ((a ? b : 13098) * (a | (14'd13851 & ((14'd6931 ^ b) ^ b))));
            
            4'd10: result_0117 = (a + ((a & 14'd1577) - 14'd8627));
            
            4'd11: result_0117 = (b | (~b));
            
            4'd12: result_0117 = ((~14'd15327) | ((((14'd14503 * 14'd11310) ^ 14'd1465) ^ (14'd13994 ? 14'd7418 : 12247)) * a));
            
            4'd13: result_0117 = (((((14'd9600 - 14'd1713) * (14'd6997 * a)) ? ((14'd3068 * b) >> 3) : 7299) & (((14'd11195 >> 2) ? (14'd11748 << 3) : 13350) << 2)) >> 3);
            
            4'd14: result_0117 = ((~((a - a) ? b : 10275)) << 2);
            
            default: result_0117 = a;
        endcase
    end

endmodule
        