
module simple_alu_0782(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0782
);

    always @(*) begin
        case(op)
            
            4'd0: result_0782 = ((b ^ a) - (((~(14'd3865 & 14'd7118)) & a) & ((14'd5338 | (b ? a : 6829)) << 3)));
            
            4'd1: result_0782 = ((((~a) | ((14'd11867 & 14'd153) ^ (a ? a : 15179))) | 14'd14506) + 14'd2047);
            
            4'd2: result_0782 = ((b & a) - (((b + (a + 14'd16128)) << 3) - (b << 3)));
            
            4'd3: result_0782 = (a ^ ((((14'd15503 ? 14'd11898 : 9644) ^ a) * 14'd10776) << 3));
            
            4'd4: result_0782 = ((14'd3890 | 14'd10380) & (~(14'd16245 * (14'd12476 >> 1))));
            
            4'd5: result_0782 = (((((b >> 3) ? 14'd12741 : 277) & 14'd9064) | (((14'd10125 | b) ? 14'd15484 : 3916) ^ 14'd13339)) ? ((~14'd1827) ^ (~((14'd15624 - 14'd2657) | (b >> 1)))) : 13049);
            
            4'd6: result_0782 = (((b ^ (~(~a))) << 3) - ((~a) - 14'd5472));
            
            4'd7: result_0782 = (~((((b << 1) - (14'd7708 >> 2)) ? b : 12208) << 2));
            
            4'd8: result_0782 = ((((14'd4890 << 2) << 1) >> 2) - 14'd1674);
            
            4'd9: result_0782 = (((((14'd8261 | 14'd2049) + 14'd7780) & (~(14'd14992 ^ 14'd9500))) ^ ((~a) + (14'd2203 * (14'd14022 >> 1)))) ? ((a ^ 14'd15529) + (((b - 14'd2426) >> 1) + ((~14'd4648) & (14'd3483 ^ 14'd8002)))) : 11192);
            
            4'd10: result_0782 = ((14'd5648 - (14'd3566 & ((a * 14'd5670) ? (b + 14'd3008) : 767))) << 2);
            
            4'd11: result_0782 = (b ^ ((~(14'd13691 << 1)) * (((14'd3975 ? 14'd4106 : 9503) | (14'd14077 * 14'd6792)) << 2)));
            
            default: result_0782 = 14'd5392;
        endcase
    end

endmodule
        