
module simple_alu_0058(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0058
);

    always @(*) begin
        case(op)
            
            4'd0: result_0058 = ((((14'd12177 & (14'd2738 * a)) << 3) << 3) << 3);
            
            4'd1: result_0058 = (b & ((b + 14'd5306) >> 1));
            
            4'd2: result_0058 = (((((14'd10875 >> 2) ^ b) * (~(~a))) >> 2) + 14'd14138);
            
            4'd3: result_0058 = (~((b * (14'd4332 + (b << 2))) >> 3));
            
            4'd4: result_0058 = ((14'd4244 + a) >> 3);
            
            4'd5: result_0058 = ((a ^ (14'd3758 * (~(a | 14'd6670)))) & ((~((~a) * (14'd3715 * 14'd826))) << 3));
            
            4'd6: result_0058 = (((b - ((14'd10403 ? b : 14181) << 1)) + (((14'd858 ? 14'd1385 : 2622) ^ (14'd14807 + b)) - ((14'd5701 ^ 14'd2312) & (14'd4794 >> 3)))) ? b : 15094);
            
            4'd7: result_0058 = (((a * ((b ? a : 3782) - (14'd2142 & b))) * 14'd3875) - (~(~b)));
            
            4'd8: result_0058 = ((~(b ^ b)) | (14'd7138 | 14'd7357));
            
            4'd9: result_0058 = (((b >> 3) * (((14'd11919 << 3) * 14'd8340) >> 2)) ^ 14'd422);
            
            4'd10: result_0058 = (14'd3183 ^ ((((a * 14'd1957) * (~14'd11803)) << 3) << 3));
            
            4'd11: result_0058 = (~((14'd695 >> 1) ? ((14'd109 - (14'd2528 ? 14'd15532 : 4444)) << 2) : 15703));
            
            4'd12: result_0058 = (b | ((14'd3354 ? 14'd10989 : 61) << 1));
            
            4'd13: result_0058 = ((14'd7407 >> 1) ^ b);
            
            default: result_0058 = a;
        endcase
    end

endmodule
        