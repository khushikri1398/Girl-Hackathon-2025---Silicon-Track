
module simple_alu_0502(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0502
);

    always @(*) begin
        case(op)
            
            4'd0: result_0502 = ((((14'd10947 * (14'd7714 ^ b)) >> 3) | (((14'd1015 ^ 14'd9442) ? (14'd5595 + 14'd8245) : 7239) | ((~b) & (~b)))) - ((b & ((b & b) ? (14'd11182 << 2) : 11563)) - (14'd13514 & ((14'd6415 ^ 14'd9205) + 14'd3137))));
            
            4'd1: result_0502 = ((b & (((~a) ? a : 11765) | ((14'd5130 >> 1) | 14'd166))) & ((((~14'd14685) ^ 14'd10201) - ((a + 14'd15586) | 14'd2116)) - 14'd14887));
            
            4'd2: result_0502 = ((14'd7044 ? ((b | (b + a)) | (b | (b | 14'd14369))) : 13522) << 1);
            
            4'd3: result_0502 = (~((((14'd2842 | a) * 14'd406) * (b & (14'd13924 + a))) - (14'd3215 | ((14'd13174 * 14'd133) & (14'd8867 | 14'd7200)))));
            
            4'd4: result_0502 = ((b + ((~14'd12584) >> 3)) ^ (14'd6352 * 14'd12711));
            
            4'd5: result_0502 = (((~14'd15574) ^ 14'd10958) ^ (((b << 2) >> 2) * ((b + (14'd7676 | 14'd7913)) ^ 14'd2846)));
            
            4'd6: result_0502 = (a << 1);
            
            4'd7: result_0502 = (14'd3973 | ((((b ? 14'd9419 : 10337) ^ (~14'd5542)) - ((14'd3995 ^ 14'd4163) - 14'd2829)) - ((14'd15590 + a) << 3)));
            
            4'd8: result_0502 = ((~(b - 14'd2611)) - (((b >> 3) + (14'd4160 ? (14'd6098 - 14'd11560) : 14332)) * (~b)));
            
            4'd9: result_0502 = ((14'd6449 ^ (((14'd12134 << 2) >> 2) | ((14'd5962 + 14'd3623) ? 14'd7876 : 1446))) >> 2);
            
            4'd10: result_0502 = ((14'd15507 & ((14'd13641 ^ (a - 14'd13526)) & ((a | 14'd11813) >> 1))) >> 2);
            
            default: result_0502 = 14'd13798;
        endcase
    end

endmodule
        