
module simple_alu_0549(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0549
);

    always @(*) begin
        case(op)
            
            4'd0: result_0549 = (14'd4873 & (14'd10150 * (((14'd13865 << 2) | (14'd3503 & 14'd8979)) * (b + (14'd11815 >> 3)))));
            
            4'd1: result_0549 = (b & ((b ? ((14'd11967 & b) - (14'd8282 - 14'd11805)) : 13332) - (14'd8674 - ((14'd8912 + 14'd5046) >> 3))));
            
            4'd2: result_0549 = ((((14'd4819 | (b << 1)) * 14'd2420) - 14'd3944) ? (((~(b << 3)) ^ 14'd9880) - (14'd8625 ? ((b - 14'd10623) >> 3) : 16074)) : 5785);
            
            4'd3: result_0549 = ((((14'd6132 >> 1) * (b * (14'd14763 * 14'd7761))) ^ (~(a ? (14'd11890 >> 2) : 15078))) + b);
            
            4'd4: result_0549 = ((b << 2) | 14'd5592);
            
            4'd5: result_0549 = ((14'd3473 & ((14'd12084 << 1) | ((14'd1489 ^ 14'd11894) | b))) + (14'd7520 + (((14'd9914 | 14'd1718) * (14'd10197 << 3)) >> 1)));
            
            4'd6: result_0549 = ((14'd10174 - (a << 3)) >> 1);
            
            4'd7: result_0549 = (a | (14'd3748 ? (14'd15210 | 14'd748) : 5810));
            
            4'd8: result_0549 = (((14'd15385 | ((b << 1) - (14'd14054 >> 3))) << 2) << 1);
            
            4'd9: result_0549 = ((~b) ^ ((((a & b) >> 2) << 2) + (14'd8737 >> 1)));
            
            4'd10: result_0549 = (14'd12221 ? b : 9578);
            
            default: result_0549 = b;
        endcase
    end

endmodule
        