
module simple_alu_0730(
    input [13:0] a, b,
    input [3:0] op,
    output reg [13:0] result_0730
);

    always @(*) begin
        case(op)
            
            4'd0: result_0730 = (((((14'd6431 + 14'd12561) - (14'd6364 ? 14'd11995 : 4323)) ? b : 5890) * ((b + (14'd4984 >> 2)) ^ ((~b) * (~14'd6072)))) | (~((14'd750 * a) << 2)));
            
            4'd1: result_0730 = ((14'd7369 ^ (a & a)) ? (b | (14'd8815 * ((14'd4850 | b) ? 14'd10155 : 5356))) : 9723);
            
            4'd2: result_0730 = ((b ^ 14'd15448) >> 2);
            
            4'd3: result_0730 = ((14'd5503 ? ((14'd10957 | (14'd2138 * 14'd8761)) | ((b & 14'd731) ? (14'd3455 ^ 14'd12579) : 8698)) : 1420) + ((((b & 14'd8015) - (14'd5424 * 14'd5858)) * 14'd4230) ^ (~((14'd3438 - a) ? (14'd7466 ? 14'd3129 : 11258) : 12316))));
            
            4'd4: result_0730 = (((14'd5202 * (b ^ (b ? a : 13119))) - (~(b ^ (14'd11337 >> 2)))) | (14'd1701 - (((14'd6261 + b) | b) << 1)));
            
            4'd5: result_0730 = (a ? ((14'd6373 << 1) + (a ^ ((14'd9307 >> 1) ^ (14'd2499 - 14'd6544)))) : 13597);
            
            4'd6: result_0730 = (14'd14056 >> 3);
            
            4'd7: result_0730 = (((14'd9801 << 1) * ((b >> 3) + ((b + a) - b))) << 1);
            
            4'd8: result_0730 = (((a - 14'd4176) - ((~(14'd13183 << 3)) + ((b ? a : 14840) & (14'd542 << 2)))) - (((a + (14'd6737 >> 1)) - (b | (b & 14'd2105))) >> 3));
            
            4'd9: result_0730 = ((((b | (~14'd12325)) - b) * (((a | 14'd13302) - (14'd8243 + 14'd6834)) ^ (~(14'd11102 | 14'd8578)))) - ((b ^ ((14'd16243 | 14'd14642) + a)) + (((a * 14'd13996) + 14'd2225) * 14'd11590)));
            
            4'd10: result_0730 = (((14'd12800 + (~(a << 3))) ^ (((~a) ? (~14'd1291) : 8275) * ((a ? 14'd3922 : 3013) ? 14'd4031 : 12342))) + 14'd5995);
            
            4'd11: result_0730 = (14'd9057 << 2);
            
            default: result_0730 = 14'd129;
        endcase
    end

endmodule
        